<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 2007" registration="Splash Software" version="DEBUG Build">
    <CONTACT name="GeoLogix AG" street="Muristrasse 60" city="Bern" zip="3006" country="CH" phone="+41 31 356 80 56" fax="+41 31 356 80 81" email="info@splash-software.ch" internet="http://www.splash-software.ch" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Nottwil" name="Schweizerische Masters Meisterschaften" name.en="Swiss Masters Championships" course="SCM" deadline="2009-09-07" nation="SUI" organizer="Schwimmverein Emmen" state="LU" timing="AUTOMATIC" type="SUI.MCS">
      <AGEDATE value="2009-09-27" type="YEAR" />
      <POOL name="Hallenbad -- Schweiz. Paraplegikerzentrum" lanemin="1" lanemax="6" />
      <POINTTABLE pointtableid="1008" name="DSV Master Performance Table" version="2004" />
      <CONTACT city="Hildisrieden" email="info@sv-emmen.ch" internet="www.sv-emmen.ch" name="Daniel Kuratli" street="Länzeweid 33b" zip="6024" />
      <SESSIONS>
        <SESSION date="2009-09-26" daytime="13:00" name="Samstag -- Einzelwettkämpfe" number="1" officialmeeting="12:15" teamleadermeeting="12:00" warmupfrom="11:30" warmupuntil="12:45">
          <EVENTS>
            <EVENT eventid="1054" daytime="13:00" gender="F" number="1" order="1" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1070" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="1056" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7170" />
                    <RANKING order="2" place="2" resultid="6964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1057" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7848" />
                    <RANKING order="2" place="2" resultid="7278" />
                    <RANKING order="3" place="3" resultid="7554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1058" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6931" />
                    <RANKING order="2" place="2" resultid="7276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1059" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1060" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1061" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7148" />
                    <RANKING order="2" place="-1" resultid="7214" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1065" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1066" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1067" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1068" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1069" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="6581" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7525" />
                    <RANKING order="2" place="2" resultid="7484" />
                    <RANKING order="3" place="3" resultid="7535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6582" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="6580" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7554" />
                    <RANKING order="2" place="2" resultid="7567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6583" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="10537" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7848" />
                    <RANKING order="2" place="2" resultid="6931" />
                    <RANKING order="3" place="3" resultid="7170" />
                    <RANKING order="4" place="4" resultid="7278" />
                    <RANKING order="5" place="5" resultid="7087" />
                    <RANKING order="6" place="6" resultid="7554" />
                    <RANKING order="7" place="7" resultid="7525" />
                    <RANKING order="8" place="8" resultid="6964" />
                    <RANKING order="9" place="9" resultid="7276" />
                    <RANKING order="10" place="10" resultid="7484" />
                    <RANKING order="11" place="11" resultid="7567" />
                    <RANKING order="12" place="12" resultid="6981" />
                    <RANKING order="13" place="13" resultid="6996" />
                    <RANKING order="14" place="14" resultid="7148" />
                    <RANKING order="15" place="15" resultid="7535" />
                    <RANKING order="16" place="-1" resultid="7214" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8535" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8536" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8537" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="13:15" gender="M" number="2" order="2" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11154" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11155" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7176" />
                    <RANKING order="2" place="2" resultid="7573" />
                    <RANKING order="3" place="-1" resultid="7151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11156" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7185" />
                    <RANKING order="2" place="-1" resultid="7499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11157" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7140" />
                    <RANKING order="2" place="2" resultid="7604" />
                    <RANKING order="3" place="-1" resultid="7093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11158" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7199" />
                    <RANKING order="2" place="2" resultid="7869" />
                    <RANKING order="3" place="3" resultid="6897" />
                    <RANKING order="4" place="4" resultid="7260" />
                    <RANKING order="5" place="5" resultid="7612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11159" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11160" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7125" />
                    <RANKING order="2" place="2" resultid="6989" />
                    <RANKING order="3" place="3" resultid="7252" />
                    <RANKING order="4" place="4" resultid="7235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11161" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6793" />
                    <RANKING order="2" place="-1" resultid="7230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11162" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7219" />
                    <RANKING order="2" place="2" resultid="6973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11163" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11164" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11165" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11166" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11167" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11168" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11169" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11170" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11171" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7612" />
                    <RANKING order="2" place="2" resultid="7604" />
                    <RANKING order="3" place="3" resultid="7511" />
                    <RANKING order="4" place="4" resultid="7573" />
                    <RANKING order="5" place="-1" resultid="7499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11172" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11173" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7199" />
                    <RANKING order="2" place="2" resultid="7176" />
                    <RANKING order="3" place="3" resultid="7869" />
                    <RANKING order="4" place="4" resultid="7140" />
                    <RANKING order="5" place="5" resultid="7185" />
                    <RANKING order="6" place="6" resultid="7125" />
                    <RANKING order="7" place="7" resultid="6793" />
                    <RANKING order="8" place="8" resultid="6897" />
                    <RANKING order="9" place="9" resultid="6989" />
                    <RANKING order="10" place="10" resultid="7260" />
                    <RANKING order="11" place="11" resultid="7252" />
                    <RANKING order="12" place="12" resultid="7612" />
                    <RANKING order="13" place="13" resultid="7235" />
                    <RANKING order="14" place="14" resultid="7219" />
                    <RANKING order="15" place="15" resultid="7511" />
                    <RANKING order="16" place="16" resultid="6973" />
                    <RANKING order="17" place="17" resultid="7296" />
                    <RANKING order="18" place="18" resultid="6828" />
                    <RANKING order="19" place="19" resultid="7604" />
                    <RANKING order="20" place="20" resultid="7573" />
                    <RANKING order="21" place="21" resultid="7599" />
                    <RANKING order="22" place="-1" resultid="7151" />
                    <RANKING order="23" place="-1" resultid="7093" />
                    <RANKING order="24" place="-1" resultid="7499" />
                    <RANKING order="25" place="-1" resultid="7230" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8538" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8539" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8540" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8541" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1282" daytime="13:35" gender="F" number="3" order="3" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11174" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6808" />
                    <RANKING order="2" place="2" resultid="6879" />
                    <RANKING order="3" place="3" resultid="7562" />
                    <RANKING order="4" place="-1" resultid="7630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11175" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11176" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11177" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11178" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11179" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11180" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11181" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11182" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11183" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11184" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11185" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11186" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11187" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11188" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11189" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7585" />
                    <RANKING order="2" place="2" resultid="7548" />
                    <RANKING order="3" place="3" resultid="7592" />
                    <RANKING order="4" place="4" resultid="7542" />
                    <RANKING order="5" place="5" resultid="7536" />
                    <RANKING order="6" place="6" resultid="7490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11190" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11191" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7556" />
                    <RANKING order="2" place="-1" resultid="7630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11192" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11193" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6808" />
                    <RANKING order="2" place="2" resultid="7001" />
                    <RANKING order="3" place="3" resultid="6879" />
                    <RANKING order="4" place="4" resultid="7114" />
                    <RANKING order="5" place="5" resultid="7585" />
                    <RANKING order="6" place="6" resultid="7556" />
                    <RANKING order="7" place="7" resultid="7300" />
                    <RANKING order="8" place="8" resultid="7166" />
                    <RANKING order="9" place="9" resultid="7163" />
                    <RANKING order="10" place="10" resultid="7548" />
                    <RANKING order="11" place="11" resultid="7562" />
                    <RANKING order="12" place="12" resultid="7592" />
                    <RANKING order="13" place="13" resultid="7542" />
                    <RANKING order="14" place="14" resultid="7536" />
                    <RANKING order="15" place="15" resultid="7490" />
                    <RANKING order="16" place="-1" resultid="7630" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8542" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8543" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8544" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1284" daytime="13:45" gender="M" number="4" order="4" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11194" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6859" />
                    <RANKING order="2" place="2" resultid="7505" />
                    <RANKING order="3" place="3" resultid="7622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11195" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7257" />
                    <RANKING order="2" place="2" resultid="6864" />
                    <RANKING order="3" place="3" resultid="7152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11196" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6819" />
                    <RANKING order="2" place="2" resultid="6947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11197" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7334" />
                    <RANKING order="2" place="2" resultid="7819" />
                    <RANKING order="3" place="-1" resultid="7879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11198" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7082" />
                    <RANKING order="2" place="2" resultid="6916" />
                    <RANKING order="3" place="3" resultid="7608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11199" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7340" />
                    <RANKING order="2" place="2" resultid="7269" />
                    <RANKING order="3" place="3" resultid="6908" />
                    <RANKING order="4" place="4" resultid="7493" />
                    <RANKING order="5" place="5" resultid="7616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11200" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6923" />
                    <RANKING order="2" place="2" resultid="6990" />
                    <RANKING order="3" place="3" resultid="7857" />
                    <RANKING order="4" place="-1" resultid="7253" />
                    <RANKING order="5" place="-1" resultid="7813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11201" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7133" />
                    <RANKING order="2" place="2" resultid="6775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11202" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11203" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11204" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11205" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11206" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11207" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11208" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11209" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11210" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11211" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7608" />
                    <RANKING order="2" place="2" resultid="7493" />
                    <RANKING order="3" place="3" resultid="7616" />
                    <RANKING order="4" place="4" resultid="7505" />
                    <RANKING order="5" place="5" resultid="7622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11212" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11213" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7334" />
                    <RANKING order="2" place="2" resultid="7340" />
                    <RANKING order="3" place="3" resultid="7819" />
                    <RANKING order="4" place="4" resultid="7257" />
                    <RANKING order="5" place="5" resultid="6819" />
                    <RANKING order="6" place="6" resultid="6864" />
                    <RANKING order="7" place="7" resultid="7133" />
                    <RANKING order="8" place="8" resultid="7082" />
                    <RANKING order="9" place="9" resultid="7269" />
                    <RANKING order="10" place="10" resultid="6916" />
                    <RANKING order="11" place="11" resultid="6859" />
                    <RANKING order="12" place="12" resultid="6923" />
                    <RANKING order="13" place="13" resultid="6775" />
                    <RANKING order="14" place="14" resultid="6947" />
                    <RANKING order="15" place="15" resultid="6990" />
                    <RANKING order="16" place="16" resultid="7220" />
                    <RANKING order="17" place="17" resultid="7152" />
                    <RANKING order="18" place="18" resultid="6781" />
                    <RANKING order="19" place="19" resultid="6908" />
                    <RANKING order="20" place="20" resultid="7857" />
                    <RANKING order="21" place="21" resultid="7608" />
                    <RANKING order="22" place="22" resultid="7666" />
                    <RANKING order="23" place="23" resultid="7493" />
                    <RANKING order="24" place="24" resultid="7505" />
                    <RANKING order="25" place="25" resultid="7671" />
                    <RANKING order="26" place="26" resultid="7616" />
                    <RANKING order="27" place="27" resultid="7622" />
                    <RANKING order="28" place="-1" resultid="7879" />
                    <RANKING order="29" place="-1" resultid="7253" />
                    <RANKING order="30" place="-1" resultid="7813" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8545" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8546" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8547" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8548" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8549" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1286" daytime="13:55" gender="F" number="5" order="5" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11214" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6868" />
                    <RANKING order="2" place="2" resultid="7569" />
                    <RANKING order="3" place="3" resultid="7579" />
                    <RANKING order="4" place="4" resultid="7581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11215" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11216" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11217" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11218" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11219" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7088" />
                    <RANKING order="2" place="2" resultid="7109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11220" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11221" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11222" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11223" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11224" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11225" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11226" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11227" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11228" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11229" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7530" />
                    <RANKING order="2" place="2" resultid="7486" />
                    <RANKING order="3" place="3" resultid="7481" />
                    <RANKING order="4" place="4" resultid="7596" />
                    <RANKING order="5" place="5" resultid="7539" />
                    <RANKING order="6" place="6" resultid="7492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11230" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11231" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7569" />
                    <RANKING order="2" place="2" resultid="7579" />
                    <RANKING order="3" place="3" resultid="7581" />
                    <RANKING order="4" place="4" resultid="7628" />
                    <RANKING order="5" place="5" resultid="7510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11232" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11233" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7088" />
                    <RANKING order="2" place="2" resultid="7109" />
                    <RANKING order="3" place="3" resultid="6868" />
                    <RANKING order="4" place="4" resultid="7530" />
                    <RANKING order="5" place="5" resultid="6982" />
                    <RANKING order="6" place="6" resultid="7103" />
                    <RANKING order="7" place="7" resultid="7486" />
                    <RANKING order="8" place="8" resultid="7569" />
                    <RANKING order="9" place="9" resultid="7481" />
                    <RANKING order="10" place="10" resultid="7596" />
                    <RANKING order="11" place="11" resultid="7579" />
                    <RANKING order="12" place="12" resultid="7581" />
                    <RANKING order="13" place="13" resultid="7628" />
                    <RANKING order="14" place="14" resultid="7539" />
                    <RANKING order="15" place="15" resultid="7492" />
                    <RANKING order="16" place="16" resultid="7510" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8550" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8551" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8552" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1288" daytime="14:10" gender="M" number="6" order="6" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11234" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11235" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7576" />
                    <RANKING order="2" place="-1" resultid="7574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11236" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6820" />
                    <RANKING order="2" place="2" resultid="7186" />
                    <RANKING order="3" place="3" resultid="7837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11237" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6845" />
                    <RANKING order="2" place="2" resultid="6906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11238" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7120" />
                    <RANKING order="2" place="2" resultid="6917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11239" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7550" />
                    <RANKING order="2" place="2" resultid="7496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11240" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6912" />
                    <RANKING order="2" place="2" resultid="7006" />
                    <RANKING order="3" place="-1" resultid="7814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11241" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11242" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11243" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11244" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11245" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11246" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11247" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11248" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11249" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7601" />
                    <RANKING order="2" place="2" resultid="7522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11250" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11251" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7550" />
                    <RANKING order="2" place="2" resultid="7496" />
                    <RANKING order="3" place="3" resultid="7576" />
                    <RANKING order="4" place="4" resultid="7624" />
                    <RANKING order="5" place="-1" resultid="7574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11252" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11253" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6845" />
                    <RANKING order="2" place="2" resultid="6820" />
                    <RANKING order="3" place="3" resultid="6906" />
                    <RANKING order="4" place="4" resultid="6912" />
                    <RANKING order="5" place="5" resultid="7186" />
                    <RANKING order="6" place="6" resultid="7837" />
                    <RANKING order="7" place="7" resultid="7120" />
                    <RANKING order="8" place="8" resultid="6917" />
                    <RANKING order="9" place="9" resultid="6974" />
                    <RANKING order="10" place="10" resultid="7550" />
                    <RANKING order="11" place="11" resultid="7006" />
                    <RANKING order="12" place="12" resultid="6786" />
                    <RANKING order="13" place="13" resultid="6829" />
                    <RANKING order="14" place="14" resultid="7496" />
                    <RANKING order="15" place="15" resultid="7576" />
                    <RANKING order="16" place="16" resultid="7601" />
                    <RANKING order="17" place="17" resultid="7522" />
                    <RANKING order="18" place="18" resultid="7672" />
                    <RANKING order="19" place="19" resultid="7624" />
                    <RANKING order="20" place="-1" resultid="7574" />
                    <RANKING order="21" place="-1" resultid="7814" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8553" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8554" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8555" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8556" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1290" daytime="14:25" gender="F" number="7" order="7" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11254" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11255" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11256" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7279" />
                    <RANKING order="2" place="2" resultid="7558" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11257" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11258" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11259" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11260" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7215" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11261" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11262" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11263" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11264" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11265" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11266" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11267" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11268" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11269" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11270" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11271" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7558" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11272" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11273" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6967" />
                    <RANKING order="2" place="2" resultid="7279" />
                    <RANKING order="3" place="3" resultid="7558" />
                    <RANKING order="4" place="4" resultid="8723" />
                    <RANKING order="5" place="-1" resultid="7215" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8557" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1292" daytime="14:25" gender="M" number="8" order="8" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11274" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11275" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6959" />
                    <RANKING order="2" place="2" resultid="7177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11276" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6948" />
                    <RANKING order="2" place="2" resultid="7187" />
                    <RANKING order="3" place="-1" resultid="7502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11277" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7880" />
                    <RANKING order="2" place="2" resultid="7606" />
                    <RANKING order="3" place="-1" resultid="7097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11278" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7870" />
                    <RANKING order="2" place="2" resultid="6898" />
                    <RANKING order="3" place="3" resultid="7613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11279" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11280" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6924" />
                    <RANKING order="2" place="2" resultid="7126" />
                    <RANKING order="3" place="3" resultid="6904" />
                    <RANKING order="4" place="4" resultid="7007" />
                    <RANKING order="5" place="5" resultid="7858" />
                    <RANKING order="6" place="6" resultid="7254" />
                    <RANKING order="7" place="7" resultid="8532" />
                    <RANKING order="8" place="8" resultid="7158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11281" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11282" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11283" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11284" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11285" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11286" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11287" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11288" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11289" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11290" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11291" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7613" />
                    <RANKING order="2" place="2" resultid="7606" />
                    <RANKING order="3" place="-1" resultid="7502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11292" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11293" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6959" />
                    <RANKING order="2" place="2" resultid="7177" />
                    <RANKING order="3" place="3" resultid="7870" />
                    <RANKING order="4" place="4" resultid="6801" />
                    <RANKING order="5" place="5" resultid="7880" />
                    <RANKING order="6" place="6" resultid="6924" />
                    <RANKING order="7" place="7" resultid="6948" />
                    <RANKING order="8" place="8" resultid="7126" />
                    <RANKING order="9" place="9" resultid="6904" />
                    <RANKING order="10" place="10" resultid="7187" />
                    <RANKING order="11" place="11" resultid="6794" />
                    <RANKING order="12" place="12" resultid="6898" />
                    <RANKING order="13" place="13" resultid="7221" />
                    <RANKING order="14" place="14" resultid="7007" />
                    <RANKING order="15" place="15" resultid="7858" />
                    <RANKING order="16" place="16" resultid="7254" />
                    <RANKING order="17" place="17" resultid="8532" />
                    <RANKING order="18" place="18" resultid="7613" />
                    <RANKING order="19" place="19" resultid="7158" />
                    <RANKING order="20" place="20" resultid="7606" />
                    <RANKING order="21" place="21" resultid="6782" />
                    <RANKING order="22" place="-1" resultid="7502" />
                    <RANKING order="23" place="-1" resultid="7097" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8558" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8559" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8560" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8561" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1294" daytime="14:35" gender="F" number="9" order="9" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11294" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6809" />
                    <RANKING order="2" place="2" resultid="6869" />
                    <RANKING order="3" place="3" resultid="7571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11295" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11296" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11297" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7272" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11298" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6968" />
                    <RANKING order="2" place="2" resultid="7115" />
                    <RANKING order="3" place="3" resultid="7104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11299" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11300" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11301" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11302" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11303" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11304" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11305" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11306" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11307" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11308" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11309" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7531" />
                    <RANKING order="2" place="2" resultid="7488" />
                    <RANKING order="3" place="3" resultid="7587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11310" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11311" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7560" />
                    <RANKING order="2" place="2" resultid="7571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11312" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11313" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7272" />
                    <RANKING order="2" place="2" resultid="6809" />
                    <RANKING order="3" place="3" resultid="7174" />
                    <RANKING order="4" place="4" resultid="6968" />
                    <RANKING order="5" place="5" resultid="7531" />
                    <RANKING order="6" place="6" resultid="7115" />
                    <RANKING order="7" place="7" resultid="6869" />
                    <RANKING order="8" place="8" resultid="7571" />
                    <RANKING order="9" place="9" resultid="7104" />
                    <RANKING order="10" place="10" resultid="7560" />
                    <RANKING order="11" place="11" resultid="6983" />
                    <RANKING order="12" place="12" resultid="7488" />
                    <RANKING order="13" place="13" resultid="7587" />
                    <RANKING order="14" place="14" resultid="7487" />
                    <RANKING order="15" place="15" resultid="6832" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8562" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8563" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8564" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1296" daytime="14:45" gender="M" number="10" order="10" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11314" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11315" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6865" />
                    <RANKING order="2" place="2" resultid="6874" />
                    <RANKING order="3" place="-1" resultid="7258" />
                    <RANKING order="4" place="-1" resultid="7577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11316" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6821" />
                    <RANKING order="2" place="2" resultid="7838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11317" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7343" />
                    <RANKING order="2" place="2" resultid="7820" />
                    <RANKING order="3" place="3" resultid="7607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11318" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6918" />
                    <RANKING order="2" place="2" resultid="6934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11319" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7551" />
                    <RANKING order="2" place="-1" resultid="7241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11320" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7255" />
                    <RANKING order="2" place="2" resultid="7008" />
                    <RANKING order="3" place="-1" resultid="6913" />
                    <RANKING order="4" place="-1" resultid="7815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11321" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11322" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11323" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11324" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6830" />
                    <RANKING order="2" place="-1" resultid="7245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11325" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11326" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11327" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11328" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11329" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11330" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11331" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7551" />
                    <RANKING order="2" place="2" resultid="7607" />
                    <RANKING order="3" place="-1" resultid="7577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11332" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11333" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7343" />
                    <RANKING order="2" place="2" resultid="7820" />
                    <RANKING order="3" place="3" resultid="6865" />
                    <RANKING order="4" place="4" resultid="6874" />
                    <RANKING order="5" place="5" resultid="6821" />
                    <RANKING order="6" place="6" resultid="6918" />
                    <RANKING order="7" place="7" resultid="7838" />
                    <RANKING order="8" place="8" resultid="7255" />
                    <RANKING order="9" place="9" resultid="7008" />
                    <RANKING order="10" place="10" resultid="6934" />
                    <RANKING order="11" place="11" resultid="7222" />
                    <RANKING order="12" place="12" resultid="6830" />
                    <RANKING order="13" place="13" resultid="7551" />
                    <RANKING order="14" place="14" resultid="7607" />
                    <RANKING order="15" place="15" resultid="6787" />
                    <RANKING order="16" place="-1" resultid="7258" />
                    <RANKING order="17" place="-1" resultid="6913" />
                    <RANKING order="18" place="-1" resultid="7815" />
                    <RANKING order="19" place="-1" resultid="7241" />
                    <RANKING order="20" place="-1" resultid="7577" />
                    <RANKING order="21" place="-1" resultid="7245" />
                    <RANKING order="22" place="-1" resultid="7134" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8565" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8566" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8567" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1298" daytime="14:55" gender="F" number="11" order="11" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11334" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6880" />
                    <RANKING order="2" place="2" resultid="6870" />
                    <RANKING order="3" place="3" resultid="7565" />
                    <RANKING order="4" place="4" resultid="7629" />
                    <RANKING order="5" place="5" resultid="7578" />
                    <RANKING order="6" place="6" resultid="7561" />
                    <RANKING order="7" place="7" resultid="7580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11335" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11336" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7849" />
                    <RANKING order="2" place="2" resultid="7552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11337" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7277" />
                    <RANKING order="2" place="2" resultid="7625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11338" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7116" />
                    <RANKING order="2" place="2" resultid="7105" />
                    <RANKING order="3" place="3" resultid="6938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11339" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11340" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7149" />
                    <RANKING order="2" place="2" resultid="7508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11341" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11342" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11343" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11344" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11345" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11346" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11347" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11348" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11349" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7523" />
                    <RANKING order="2" place="2" resultid="7482" />
                    <RANKING order="3" place="3" resultid="7582" />
                    <RANKING order="4" place="4" resultid="7545" />
                    <RANKING order="5" place="5" resultid="7590" />
                    <RANKING order="6" place="6" resultid="7533" />
                    <RANKING order="7" place="7" resultid="7489" />
                    <RANKING order="8" place="-1" resultid="7540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11350" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11351" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7552" />
                    <RANKING order="2" place="2" resultid="7565" />
                    <RANKING order="3" place="3" resultid="7578" />
                    <RANKING order="4" place="4" resultid="7629" />
                    <RANKING order="5" place="5" resultid="7580" />
                    <RANKING order="6" place="6" resultid="7625" />
                    <RANKING order="7" place="7" resultid="7508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11352" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11353" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7277" />
                    <RANKING order="2" place="2" resultid="7002" />
                    <RANKING order="3" place="3" resultid="7849" />
                    <RANKING order="4" place="4" resultid="7552" />
                    <RANKING order="5" place="5" resultid="7523" />
                    <RANKING order="6" place="6" resultid="6880" />
                    <RANKING order="7" place="6" resultid="6965" />
                    <RANKING order="8" place="8" resultid="6870" />
                    <RANKING order="9" place="9" resultid="7565" />
                    <RANKING order="10" place="10" resultid="7116" />
                    <RANKING order="11" place="11" resultid="7105" />
                    <RANKING order="12" place="12" resultid="7482" />
                    <RANKING order="13" place="13" resultid="7301" />
                    <RANKING order="14" place="14" resultid="7582" />
                    <RANKING order="15" place="15" resultid="6938" />
                    <RANKING order="16" place="16" resultid="7149" />
                    <RANKING order="17" place="17" resultid="7545" />
                    <RANKING order="18" place="18" resultid="7629" />
                    <RANKING order="19" place="19" resultid="7578" />
                    <RANKING order="20" place="20" resultid="7590" />
                    <RANKING order="21" place="21" resultid="7561" />
                    <RANKING order="22" place="22" resultid="7580" />
                    <RANKING order="23" place="23" resultid="7625" />
                    <RANKING order="24" place="24" resultid="7508" />
                    <RANKING order="25" place="25" resultid="7533" />
                    <RANKING order="26" place="26" resultid="7489" />
                    <RANKING order="27" place="-1" resultid="7164" />
                    <RANKING order="28" place="-1" resultid="7540" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8569" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8570" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8571" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8572" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8573" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1300" daytime="15:10" gender="M" number="12" order="12" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11354" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6860" />
                    <RANKING order="2" place="2" resultid="7503" />
                    <RANKING order="3" place="3" resultid="7620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11355" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7178" />
                    <RANKING order="2" place="2" resultid="6960" />
                    <RANKING order="3" place="3" resultid="7259" />
                    <RANKING order="4" place="4" resultid="6875" />
                    <RANKING order="5" place="5" resultid="6841" />
                    <RANKING order="6" place="6" resultid="6886" />
                    <RANKING order="7" place="7" resultid="7575" />
                    <RANKING order="8" place="-1" resultid="7572" />
                    <RANKING order="9" place="-1" resultid="7153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11356" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6822" />
                    <RANKING order="2" place="2" resultid="6949" />
                    <RANKING order="3" place="3" resultid="7188" />
                    <RANKING order="4" place="-1" resultid="7497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11357" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6846" />
                    <RANKING order="2" place="2" resultid="6907" />
                    <RANKING order="3" place="3" resultid="7602" />
                    <RANKING order="4" place="4" resultid="7614" />
                    <RANKING order="5" place="-1" resultid="7094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11358" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7871" />
                    <RANKING order="2" place="2" resultid="6899" />
                    <RANKING order="3" place="3" resultid="7261" />
                    <RANKING order="4" place="4" resultid="7083" />
                    <RANKING order="5" place="5" resultid="7121" />
                    <RANKING order="6" place="6" resultid="6919" />
                    <RANKING order="7" place="7" resultid="7610" />
                    <RANKING order="8" place="8" resultid="8656" />
                    <RANKING order="9" place="9" resultid="6940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11359" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6802" />
                    <RANKING order="2" place="2" resultid="6909" />
                    <RANKING order="3" place="3" resultid="7618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11360" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6939" />
                    <RANKING order="2" place="2" resultid="6914" />
                    <RANKING order="3" place="3" resultid="6903" />
                    <RANKING order="4" place="4" resultid="7127" />
                    <RANKING order="5" place="5" resultid="6925" />
                    <RANKING order="6" place="6" resultid="6991" />
                    <RANKING order="7" place="7" resultid="7855" />
                    <RANKING order="8" place="8" resultid="7256" />
                    <RANKING order="9" place="9" resultid="7009" />
                    <RANKING order="10" place="10" resultid="8531" />
                    <RANKING order="11" place="11" resultid="7159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11361" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11362" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7223" />
                    <RANKING order="2" place="2" resultid="6975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11363" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11364" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11365" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11366" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11367" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11368" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11369" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7519" />
                    <RANKING order="2" place="2" resultid="7597" />
                    <RANKING order="3" place="3" resultid="7588" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11370" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11371" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7610" />
                    <RANKING order="2" place="2" resultid="7602" />
                    <RANKING order="3" place="3" resultid="8528" />
                    <RANKING order="4" place="4" resultid="7575" />
                    <RANKING order="5" place="5" resultid="7614" />
                    <RANKING order="6" place="6" resultid="7620" />
                    <RANKING order="7" place="7" resultid="7618" />
                    <RANKING order="8" place="8" resultid="7503" />
                    <RANKING order="9" place="-1" resultid="7572" />
                    <RANKING order="10" place="-1" resultid="7497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11372" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11373" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7178" />
                    <RANKING order="2" place="2" resultid="6960" />
                    <RANKING order="3" place="3" resultid="6846" />
                    <RANKING order="4" place="4" resultid="7871" />
                    <RANKING order="5" place="5" resultid="6860" />
                    <RANKING order="6" place="6" resultid="6802" />
                    <RANKING order="7" place="7" resultid="7259" />
                    <RANKING order="8" place="8" resultid="6907" />
                    <RANKING order="9" place="9" resultid="6875" />
                    <RANKING order="10" place="10" resultid="6822" />
                    <RANKING order="11" place="11" resultid="6899" />
                    <RANKING order="12" place="12" resultid="6939" />
                    <RANKING order="13" place="13" resultid="7261" />
                    <RANKING order="14" place="14" resultid="6914" />
                    <RANKING order="15" place="15" resultid="6841" />
                    <RANKING order="16" place="16" resultid="7083" />
                    <RANKING order="17" place="17" resultid="6903" />
                    <RANKING order="18" place="18" resultid="7127" />
                    <RANKING order="19" place="18" resultid="7121" />
                    <RANKING order="20" place="20" resultid="6925" />
                    <RANKING order="21" place="21" resultid="6949" />
                    <RANKING order="22" place="22" resultid="6919" />
                    <RANKING order="23" place="23" resultid="7223" />
                    <RANKING order="24" place="24" resultid="6991" />
                    <RANKING order="25" place="25" resultid="7188" />
                    <RANKING order="26" place="26" resultid="7855" />
                    <RANKING order="27" place="27" resultid="7256" />
                    <RANKING order="28" place="28" resultid="7610" />
                    <RANKING order="29" place="29" resultid="7009" />
                    <RANKING order="30" place="30" resultid="8531" />
                    <RANKING order="31" place="31" resultid="8656" />
                    <RANKING order="32" place="32" resultid="6975" />
                    <RANKING order="33" place="33" resultid="7159" />
                    <RANKING order="34" place="34" resultid="6909" />
                    <RANKING order="35" place="35" resultid="6886" />
                    <RANKING order="36" place="36" resultid="6940" />
                    <RANKING order="37" place="37" resultid="7602" />
                    <RANKING order="38" place="38" resultid="8528" />
                    <RANKING order="39" place="39" resultid="7575" />
                    <RANKING order="40" place="40" resultid="7614" />
                    <RANKING order="41" place="41" resultid="7519" />
                    <RANKING order="42" place="42" resultid="7597" />
                    <RANKING order="43" place="43" resultid="7503" />
                    <RANKING order="44" place="44" resultid="7618" />
                    <RANKING order="45" place="45" resultid="7589" />
                    <RANKING order="46" place="46" resultid="7620" />
                    <RANKING order="47" place="47" resultid="7588" />
                    <RANKING order="48" place="-1" resultid="7572" />
                    <RANKING order="49" place="-1" resultid="7497" />
                    <RANKING order="50" place="-1" resultid="7094" />
                    <RANKING order="51" place="-1" resultid="7153" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8574" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8575" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8576" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8577" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8578" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8579" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8580" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8581" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9290" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1302" daytime="15:25" gender="F" number="13" order="13" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11374" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11375" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11376" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11377" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11378" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11379" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11380" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7167" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11381" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11382" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11383" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6833" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11384" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11385" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11386" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11387" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11388" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11389" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11390" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11391" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11392" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11393" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6810" />
                    <RANKING order="2" place="2" resultid="6997" />
                    <RANKING order="3" place="3" resultid="7167" />
                    <RANKING order="4" place="4" resultid="6833" />
                    <RANKING order="5" place="5" resultid="7594" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8582" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1304" daytime="15:35" gender="M" number="14" order="14" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11394" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11395" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11396" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11397" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11398" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11399" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7270" />
                    <RANKING order="2" place="-1" resultid="7242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11400" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11401" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7135" />
                    <RANKING order="2" place="2" resultid="6776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11402" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11403" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11404" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6783" />
                    <RANKING order="2" place="2" resultid="6831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11405" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11406" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11407" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11408" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11409" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11410" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11411" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11412" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11413" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7821" />
                    <RANKING order="2" place="2" resultid="7135" />
                    <RANKING order="3" place="3" resultid="7270" />
                    <RANKING order="4" place="4" resultid="6776" />
                    <RANKING order="5" place="5" resultid="7224" />
                    <RANKING order="6" place="6" resultid="6783" />
                    <RANKING order="7" place="7" resultid="6831" />
                    <RANKING order="8" place="8" resultid="7667" />
                    <RANKING order="9" place="-1" resultid="7250" />
                    <RANKING order="10" place="-1" resultid="7154" />
                    <RANKING order="11" place="-1" resultid="7242" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8583" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8584" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-26" daytime="15:50" name="Samstag -- Staffeln" number="2">
          <EVENTS>
            <EVENT eventid="1175" daytime="15:50" gender="X" number="15" order="8" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="2000" />
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1176" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7434" />
                    <RANKING order="2" place="2" resultid="7012" />
                    <RANKING order="3" place="3" resultid="6882" />
                    <RANKING order="4" place="4" resultid="7292" />
                    <RANKING order="5" place="5" resultid="7437" />
                    <RANKING order="6" place="6" resultid="7436" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8585" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-26" daytime="16:00" name="Samstag -- 800 m" number="3">
          <EVENTS>
            <EVENT eventid="1177" daytime="16:00" gender="F" number="16" order="8" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11414" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11415" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7171" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11416" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11417" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11418" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11419" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11420" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11421" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11422" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11423" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11424" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11425" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11426" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11427" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11428" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11429" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11430" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11431" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11432" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11433" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7171" />
                    <RANKING order="2" place="2" resultid="6932" />
                    <RANKING order="3" place="3" resultid="7850" />
                    <RANKING order="4" place="4" resultid="7110" />
                    <RANKING order="5" place="5" resultid="6969" />
                    <RANKING order="6" place="6" resultid="6984" />
                    <RANKING order="7" place="7" resultid="9734" />
                    <RANKING order="8" place="8" resultid="6834" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8587" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8588" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1196" daytime="16:35" gender="M" number="17" order="9" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11434" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11435" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11436" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11437" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11438" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9741" />
                    <RANKING order="2" place="2" resultid="8750" />
                    <RANKING order="3" place="3" resultid="7262" />
                    <RANKING order="4" place="4" resultid="6935" />
                    <RANKING order="5" place="-1" resultid="7266" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11439" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11440" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7128" />
                    <RANKING order="2" place="2" resultid="6992" />
                    <RANKING order="3" place="3" resultid="9740" />
                    <RANKING order="4" place="4" resultid="7010" />
                    <RANKING order="5" place="5" resultid="9743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11441" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6795" />
                    <RANKING order="2" place="-1" resultid="7231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11442" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11443" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11444" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11445" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11446" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11447" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11448" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11449" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11450" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11451" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7513" />
                    <RANKING order="2" place="-1" resultid="7501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11452" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11453" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9741" />
                    <RANKING order="2" place="2" resultid="7141" />
                    <RANKING order="3" place="3" resultid="8750" />
                    <RANKING order="4" place="4" resultid="6795" />
                    <RANKING order="5" place="5" resultid="7128" />
                    <RANKING order="6" place="6" resultid="7262" />
                    <RANKING order="7" place="7" resultid="6992" />
                    <RANKING order="8" place="8" resultid="6976" />
                    <RANKING order="9" place="9" resultid="6935" />
                    <RANKING order="10" place="10" resultid="9740" />
                    <RANKING order="11" place="11" resultid="7010" />
                    <RANKING order="12" place="12" resultid="7297" />
                    <RANKING order="13" place="13" resultid="9743" />
                    <RANKING order="14" place="14" resultid="7513" />
                    <RANKING order="15" place="-1" resultid="7266" />
                    <RANKING order="16" place="-1" resultid="7246" />
                    <RANKING order="17" place="-1" resultid="7501" />
                    <RANKING order="18" place="-1" resultid="7231" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8589" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8590" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9736" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-27" name="Samstag  -- 1500m" number="4">
          <EVENTS>
            <EVENT eventid="7347" number="18" order="2" preveventid="-1" round="TIM">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7348" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7430" />
                    <RANKING order="2" place="2" resultid="7431" />
                    <RANKING order="3" place="3" resultid="8634" />
                    <RANKING order="4" place="4" resultid="8684" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8592" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-27" daytime="09:00" name="Sonntag -- Einzelwettkämpfe" number="7" officialmeeting="08:30" teamleadermeeting="08:15" warmupfrom="08:00" warmupuntil="08:45">
          <EVENTS>
            <EVENT eventid="1072" daytime="09:00" gender="F" number="19" order="2" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11454" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6815" />
                    <RANKING order="2" place="2" resultid="6811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11455" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7172" />
                    <RANKING order="2" place="2" resultid="7013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11456" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7851" />
                    <RANKING order="2" place="2" resultid="7280" />
                    <RANKING order="3" place="3" resultid="7555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11457" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11458" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11459" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7111" />
                    <RANKING order="2" place="-1" resultid="7089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11460" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11461" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11462" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11463" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11464" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11465" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11466" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11467" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11468" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11469" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7526" />
                    <RANKING order="2" place="2" resultid="7485" />
                    <RANKING order="3" place="3" resultid="7584" />
                    <RANKING order="4" place="4" resultid="7547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11470" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11471" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11472" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11473" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7172" />
                    <RANKING order="2" place="2" resultid="6933" />
                    <RANKING order="3" place="3" resultid="7851" />
                    <RANKING order="4" place="4" resultid="6815" />
                    <RANKING order="5" place="5" resultid="7280" />
                    <RANKING order="6" place="6" resultid="6811" />
                    <RANKING order="7" place="7" resultid="7526" />
                    <RANKING order="8" place="8" resultid="7555" />
                    <RANKING order="9" place="9" resultid="7111" />
                    <RANKING order="10" place="10" resultid="7013" />
                    <RANKING order="11" place="11" resultid="7485" />
                    <RANKING order="12" place="12" resultid="6985" />
                    <RANKING order="13" place="13" resultid="7584" />
                    <RANKING order="14" place="14" resultid="7547" />
                    <RANKING order="15" place="-1" resultid="7216" />
                    <RANKING order="16" place="-1" resultid="7089" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8593" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8594" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8595" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1157" daytime="09:25" gender="M" number="20" order="3" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11474" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11475" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11476" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6950" />
                    <RANKING order="2" place="-1" resultid="7500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11477" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7142" />
                    <RANKING order="2" place="2" resultid="7605" />
                    <RANKING order="3" place="-1" resultid="7095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11478" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7267" />
                    <RANKING order="2" place="2" resultid="7084" />
                    <RANKING order="3" place="3" resultid="6900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11479" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7512" />
                    <RANKING order="2" place="-1" resultid="7662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11480" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11481" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6796" />
                    <RANKING order="2" place="2" resultid="6922" />
                    <RANKING order="3" place="-1" resultid="7232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11482" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6977" />
                    <RANKING order="2" place="2" resultid="7225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11483" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11484" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11485" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11486" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11487" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11488" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11489" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11490" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11491" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7605" />
                    <RANKING order="2" place="2" resultid="7512" />
                    <RANKING order="3" place="-1" resultid="7500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11492" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11493" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7267" />
                    <RANKING order="2" place="2" resultid="7142" />
                    <RANKING order="3" place="3" resultid="7084" />
                    <RANKING order="4" place="4" resultid="6796" />
                    <RANKING order="5" place="5" resultid="6950" />
                    <RANKING order="6" place="6" resultid="6900" />
                    <RANKING order="7" place="7" resultid="6993" />
                    <RANKING order="8" place="8" resultid="6977" />
                    <RANKING order="9" place="9" resultid="7225" />
                    <RANKING order="10" place="10" resultid="7512" />
                    <RANKING order="11" place="11" resultid="7605" />
                    <RANKING order="12" place="12" resultid="6922" />
                    <RANKING order="13" place="-1" resultid="7662" />
                    <RANKING order="14" place="-1" resultid="7095" />
                    <RANKING order="15" place="-1" resultid="7500" />
                    <RANKING order="16" place="-1" resultid="7232" />
                    <RANKING order="17" place="-1" resultid="7247" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8596" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8597" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8598" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" daytime="09:55" gender="F" number="21" order="4" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10902" agemax="17" agemin="-1" />
                <AGEGROUP agegroupid="10903" agemax="24" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6816" />
                    <RANKING order="2" place="2" resultid="7528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10904" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="10905" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7281" />
                    <RANKING order="2" place="2" resultid="7559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10906" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10907" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10908" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="10909" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10910" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="10911" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="10912" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10913" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10914" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10915" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="10916" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="10917" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="10918" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10919" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="10920" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10921" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="10922" agemax="-1" agemin="-1" name="Klassierung nach Zeit" type="MASTERS">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7273" />
                    <RANKING order="2" place="2" resultid="6816" />
                    <RANKING order="3" place="3" resultid="7281" />
                    <RANKING order="4" place="4" resultid="6970" />
                    <RANKING order="5" place="5" resultid="7528" />
                    <RANKING order="6" place="6" resultid="7559" />
                    <RANKING order="7" place="-1" resultid="7217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11494" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7273" />
                    <RANKING order="2" place="2" resultid="6816" />
                    <RANKING order="3" place="3" resultid="7281" />
                    <RANKING order="4" place="4" resultid="6970" />
                    <RANKING order="5" place="5" resultid="7528" />
                    <RANKING order="6" place="6" resultid="7559" />
                    <RANKING order="7" place="-1" resultid="7217" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8599" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1342" daytime="10:00" gender="M" number="22" order="5" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11495" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11496" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6961" />
                    <RANKING order="2" place="2" resultid="7179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11497" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11498" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11499" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11500" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6956" />
                    <RANKING order="2" place="2" resultid="6803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11501" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7129" />
                    <RANKING order="2" place="2" resultid="7239" />
                    <RANKING order="3" place="3" resultid="7856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11502" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11503" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11504" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11505" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6784" />
                    <RANKING order="2" place="-1" resultid="7248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11506" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11507" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11508" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11509" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11510" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11511" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11512" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11513" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11514" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6961" />
                    <RANKING order="2" place="2" resultid="6956" />
                    <RANKING order="3" place="3" resultid="6803" />
                    <RANKING order="4" place="4" resultid="7179" />
                    <RANKING order="5" place="5" resultid="7196" />
                    <RANKING order="6" place="6" resultid="7129" />
                    <RANKING order="7" place="7" resultid="7226" />
                    <RANKING order="8" place="8" resultid="7239" />
                    <RANKING order="9" place="9" resultid="7856" />
                    <RANKING order="10" place="10" resultid="6784" />
                    <RANKING order="11" place="-1" resultid="7248" />
                    <RANKING order="12" place="-1" resultid="7233" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8600" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8601" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1360" daytime="10:10" gender="F" number="23" order="6" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11515" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6871" />
                    <RANKING order="2" place="2" resultid="7568" />
                    <RANKING order="3" place="3" resultid="7564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11516" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11517" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11518" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7274" />
                    <RANKING order="2" place="2" resultid="7627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11519" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11520" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11521" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11522" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11523" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11524" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11525" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11526" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11527" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11528" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11529" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11530" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7529" />
                    <RANKING order="2" place="2" resultid="9856" />
                    <RANKING order="3" place="3" resultid="7480" />
                    <RANKING order="4" place="4" resultid="7595" />
                    <RANKING order="5" place="5" resultid="7544" />
                    <RANKING order="6" place="6" resultid="7491" />
                    <RANKING order="7" place="7" resultid="7538" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11531" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11532" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7568" />
                    <RANKING order="2" place="2" resultid="7627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11533" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11534" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7274" />
                    <RANKING order="2" place="2" resultid="7529" />
                    <RANKING order="3" place="3" resultid="6871" />
                    <RANKING order="4" place="4" resultid="7568" />
                    <RANKING order="5" place="5" resultid="7106" />
                    <RANKING order="6" place="6" resultid="9856" />
                    <RANKING order="7" place="7" resultid="6986" />
                    <RANKING order="8" place="8" resultid="7480" />
                    <RANKING order="9" place="9" resultid="7595" />
                    <RANKING order="10" place="10" resultid="7564" />
                    <RANKING order="11" place="11" resultid="7627" />
                    <RANKING order="12" place="12" resultid="7544" />
                    <RANKING order="13" place="13" resultid="7491" />
                    <RANKING order="14" place="14" resultid="7538" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8602" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8603" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8604" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1378" daytime="10:20" gender="M" number="24" order="7" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11535" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7507" />
                    <RANKING order="2" place="2" resultid="7623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11536" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6876" />
                    <RANKING order="2" place="2" resultid="6842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11537" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11538" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="6847" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11539" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7876" />
                    <RANKING order="2" place="2" resultid="7122" />
                    <RANKING order="3" place="3" resultid="6920" />
                    <RANKING order="4" place="4" resultid="6901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11540" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6957" />
                    <RANKING order="2" place="2" resultid="7514" />
                    <RANKING order="3" place="3" resultid="7495" />
                    <RANKING order="4" place="4" resultid="7619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11541" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6915" />
                    <RANKING order="2" place="2" resultid="6905" />
                    <RANKING order="3" place="3" resultid="7160" />
                    <RANKING order="4" place="-1" resultid="7816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11542" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11543" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11544" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11545" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11546" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11547" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11548" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11549" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11550" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7600" />
                    <RANKING order="2" place="2" resultid="7520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11551" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11552" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7514" />
                    <RANKING order="2" place="2" resultid="7495" />
                    <RANKING order="3" place="3" resultid="7623" />
                    <RANKING order="4" place="4" resultid="7619" />
                    <RANKING order="5" place="5" resultid="7507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11553" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11554" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6957" />
                    <RANKING order="2" place="2" resultid="7876" />
                    <RANKING order="3" place="3" resultid="6876" />
                    <RANKING order="4" place="4" resultid="6915" />
                    <RANKING order="5" place="5" resultid="6842" />
                    <RANKING order="6" place="6" resultid="7839" />
                    <RANKING order="7" place="7" resultid="6905" />
                    <RANKING order="8" place="8" resultid="7122" />
                    <RANKING order="9" place="9" resultid="6978" />
                    <RANKING order="10" place="9" resultid="6920" />
                    <RANKING order="11" place="11" resultid="6901" />
                    <RANKING order="12" place="12" resultid="7514" />
                    <RANKING order="13" place="13" resultid="7160" />
                    <RANKING order="14" place="14" resultid="6788" />
                    <RANKING order="15" place="15" resultid="7495" />
                    <RANKING order="16" place="16" resultid="7600" />
                    <RANKING order="17" place="17" resultid="7520" />
                    <RANKING order="18" place="18" resultid="7673" />
                    <RANKING order="19" place="19" resultid="7507" />
                    <RANKING order="20" place="20" resultid="7619" />
                    <RANKING order="21" place="21" resultid="7623" />
                    <RANKING order="22" place="-1" resultid="7816" />
                    <RANKING order="23" place="-1" resultid="6847" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8605" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8606" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8607" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8608" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1396" daytime="10:30" gender="F" number="25" order="8" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11555" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6812" />
                    <RANKING order="2" place="2" resultid="6881" />
                    <RANKING order="3" place="-1" resultid="7563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11556" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11557" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11558" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11559" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6837" />
                    <RANKING order="2" place="2" resultid="7117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11560" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11561" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11562" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11563" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11564" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11565" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11566" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11567" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11568" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11569" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11570" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7586" />
                    <RANKING order="2" place="2" resultid="7527" />
                    <RANKING order="3" place="3" resultid="7549" />
                    <RANKING order="4" place="4" resultid="7593" />
                    <RANKING order="5" place="5" resultid="7543" />
                    <RANKING order="6" place="6" resultid="7537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11571" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11572" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11573" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11574" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6837" />
                    <RANKING order="2" place="2" resultid="6812" />
                    <RANKING order="3" place="3" resultid="7003" />
                    <RANKING order="4" place="4" resultid="7117" />
                    <RANKING order="5" place="5" resultid="6881" />
                    <RANKING order="6" place="6" resultid="7289" />
                    <RANKING order="7" place="7" resultid="7586" />
                    <RANKING order="8" place="8" resultid="7527" />
                    <RANKING order="9" place="9" resultid="6999" />
                    <RANKING order="10" place="10" resultid="7549" />
                    <RANKING order="11" place="11" resultid="7593" />
                    <RANKING order="12" place="12" resultid="7543" />
                    <RANKING order="13" place="13" resultid="7537" />
                    <RANKING order="14" place="-1" resultid="7563" />
                    <RANKING order="15" place="-1" resultid="7557" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8609" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8610" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8611" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1414" daytime="10:40" gender="M" number="26" order="9" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11575" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6861" />
                    <RANKING order="2" place="2" resultid="7506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11576" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6866" />
                    <RANKING order="2" place="-1" resultid="6852" />
                    <RANKING order="3" place="-1" resultid="7155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11577" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11578" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7822" />
                    <RANKING order="2" place="2" resultid="6943" />
                    <RANKING order="3" place="-1" resultid="7335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11579" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7085" />
                    <RANKING order="2" place="2" resultid="6921" />
                    <RANKING order="3" place="3" resultid="7609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11580" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6910" />
                    <RANKING order="2" place="2" resultid="7494" />
                    <RANKING order="3" place="3" resultid="7615" />
                    <RANKING order="4" place="-1" resultid="7341" />
                    <RANKING order="5" place="-1" resultid="7243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11581" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11582" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7136" />
                    <RANKING order="2" place="2" resultid="6777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11583" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11584" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6789" />
                    <RANKING order="2" place="2" resultid="7668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11585" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11586" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11587" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11588" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11589" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11590" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11591" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11592" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7609" />
                    <RANKING order="2" place="2" resultid="7494" />
                    <RANKING order="3" place="3" resultid="7615" />
                    <RANKING order="4" place="4" resultid="7506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11593" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11594" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7822" />
                    <RANKING order="2" place="2" resultid="7136" />
                    <RANKING order="3" place="3" resultid="6866" />
                    <RANKING order="4" place="4" resultid="6943" />
                    <RANKING order="5" place="5" resultid="7085" />
                    <RANKING order="6" place="6" resultid="6921" />
                    <RANKING order="7" place="7" resultid="6861" />
                    <RANKING order="8" place="8" resultid="6777" />
                    <RANKING order="9" place="9" resultid="7609" />
                    <RANKING order="10" place="10" resultid="7227" />
                    <RANKING order="11" place="11" resultid="6785" />
                    <RANKING order="12" place="12" resultid="6910" />
                    <RANKING order="13" place="13" resultid="6789" />
                    <RANKING order="14" place="14" resultid="7668" />
                    <RANKING order="15" place="15" resultid="7494" />
                    <RANKING order="16" place="16" resultid="7506" />
                    <RANKING order="17" place="17" resultid="7615" />
                    <RANKING order="18" place="-1" resultid="7341" />
                    <RANKING order="19" place="-1" resultid="7335" />
                    <RANKING order="20" place="-1" resultid="7155" />
                    <RANKING order="21" place="-1" resultid="6852" />
                    <RANKING order="22" place="-1" resultid="7243" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8612" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8613" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8614" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8615" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1432" daytime="10:55" gender="F" number="27" order="10" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11595" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7566" />
                    <RANKING order="2" place="2" resultid="6872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11596" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7173" />
                    <RANKING order="2" place="2" resultid="7014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11597" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7852" />
                    <RANKING order="2" place="2" resultid="7282" />
                    <RANKING order="3" place="3" resultid="7553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11598" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11599" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11600" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7112" />
                    <RANKING order="2" place="-1" resultid="7090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11601" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7290" />
                    <RANKING order="2" place="2" resultid="7509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11602" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11603" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11604" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11605" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11606" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11607" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11608" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11609" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11610" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7524" />
                    <RANKING order="2" place="2" resultid="7483" />
                    <RANKING order="3" place="3" resultid="7583" />
                    <RANKING order="4" place="4" resultid="7546" />
                    <RANKING order="5" place="5" resultid="7591" />
                    <RANKING order="6" place="6" resultid="7541" />
                    <RANKING order="7" place="7" resultid="7534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11611" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11612" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7553" />
                    <RANKING order="2" place="2" resultid="7566" />
                    <RANKING order="3" place="3" resultid="7509" />
                    <RANKING order="4" place="-1" resultid="7626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11613" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11614" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7852" />
                    <RANKING order="2" place="2" resultid="7173" />
                    <RANKING order="3" place="3" resultid="7282" />
                    <RANKING order="4" place="4" resultid="7524" />
                    <RANKING order="5" place="5" resultid="7112" />
                    <RANKING order="6" place="6" resultid="7118" />
                    <RANKING order="7" place="7" resultid="7553" />
                    <RANKING order="8" place="8" resultid="7014" />
                    <RANKING order="9" place="9" resultid="7566" />
                    <RANKING order="10" place="10" resultid="6872" />
                    <RANKING order="11" place="11" resultid="7483" />
                    <RANKING order="12" place="12" resultid="7290" />
                    <RANKING order="13" place="13" resultid="7583" />
                    <RANKING order="14" place="14" resultid="7546" />
                    <RANKING order="15" place="15" resultid="7591" />
                    <RANKING order="16" place="16" resultid="7541" />
                    <RANKING order="17" place="17" resultid="7509" />
                    <RANKING order="18" place="18" resultid="7534" />
                    <RANKING order="19" place="-1" resultid="7626" />
                    <RANKING order="20" place="-1" resultid="7004" />
                    <RANKING order="21" place="-1" resultid="7090" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8616" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8617" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8618" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8619" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1450" daytime="11:10" gender="M" number="28" order="11" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11615" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6862" />
                    <RANKING order="2" place="2" resultid="7504" />
                    <RANKING order="3" place="3" resultid="7621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11616" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6962" />
                    <RANKING order="2" place="2" resultid="7180" />
                    <RANKING order="3" place="3" resultid="6877" />
                    <RANKING order="4" place="4" resultid="6843" />
                    <RANKING order="5" place="-1" resultid="7156" />
                    <RANKING order="6" place="-1" resultid="6853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11617" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6951" />
                    <RANKING order="2" place="-1" resultid="7498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11618" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7603" />
                    <RANKING order="2" place="-1" resultid="7096" />
                    <RANKING order="3" place="-1" resultid="6848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11619" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7877" />
                    <RANKING order="2" place="2" resultid="6902" />
                    <RANKING order="3" place="3" resultid="7182" />
                    <RANKING order="4" place="4" resultid="7197" />
                    <RANKING order="5" place="5" resultid="6936" />
                    <RANKING order="6" place="6" resultid="7611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11620" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6911" />
                    <RANKING order="2" place="2" resultid="7617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11621" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7130" />
                    <RANKING order="2" place="2" resultid="6994" />
                    <RANKING order="3" place="3" resultid="7161" />
                    <RANKING order="4" place="-1" resultid="8533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11622" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6797" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11623" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11624" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11625" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11626" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11627" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11628" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11629" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11630" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7598" />
                    <RANKING order="2" place="2" resultid="7521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11631" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11632" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7611" />
                    <RANKING order="2" place="2" resultid="7603" />
                    <RANKING order="3" place="3" resultid="7621" />
                    <RANKING order="4" place="4" resultid="7617" />
                    <RANKING order="5" place="5" resultid="7504" />
                    <RANKING order="6" place="-1" resultid="7498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11633" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11634" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6962" />
                    <RANKING order="2" place="2" resultid="7180" />
                    <RANKING order="3" place="3" resultid="7877" />
                    <RANKING order="4" place="4" resultid="6877" />
                    <RANKING order="5" place="5" resultid="6862" />
                    <RANKING order="6" place="6" resultid="6902" />
                    <RANKING order="7" place="7" resultid="6843" />
                    <RANKING order="8" place="8" resultid="7182" />
                    <RANKING order="9" place="9" resultid="6797" />
                    <RANKING order="10" place="10" resultid="7197" />
                    <RANKING order="11" place="11" resultid="7130" />
                    <RANKING order="12" place="12" resultid="6951" />
                    <RANKING order="13" place="13" resultid="6994" />
                    <RANKING order="14" place="14" resultid="6936" />
                    <RANKING order="15" place="15" resultid="7611" />
                    <RANKING order="16" place="16" resultid="7228" />
                    <RANKING order="17" place="17" resultid="7161" />
                    <RANKING order="18" place="18" resultid="7603" />
                    <RANKING order="19" place="19" resultid="6911" />
                    <RANKING order="20" place="20" resultid="7521" />
                    <RANKING order="21" place="21" resultid="7598" />
                    <RANKING order="22" place="22" resultid="7617" />
                    <RANKING order="23" place="23" resultid="7504" />
                    <RANKING order="24" place="24" resultid="7621" />
                    <RANKING order="25" place="-1" resultid="8533" />
                    <RANKING order="26" place="-1" resultid="7156" />
                    <RANKING order="27" place="-1" resultid="7498" />
                    <RANKING order="28" place="-1" resultid="7096" />
                    <RANKING order="29" place="-1" resultid="6848" />
                    <RANKING order="30" place="-1" resultid="6853" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8620" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8621" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8622" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8623" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8624" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1468" daytime="11:25" gender="F" number="29" order="12" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11635" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11636" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11637" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11638" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11639" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11640" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11641" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11642" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11643" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11644" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11645" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11646" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11647" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11648" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11649" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11650" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11651" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11652" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11653" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11654" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7107" />
                    <RANKING order="2" place="2" resultid="6987" />
                    <RANKING order="3" place="3" resultid="7570" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8625" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1486" daytime="11:30" gender="M" number="30" order="13" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11655" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11656" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11657" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11658" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11659" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11660" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7271" />
                    <RANKING order="2" place="2" resultid="9092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11661" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11662" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11663" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11664" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11665" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11666" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11667" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11668" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11669" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11670" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11671" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11672" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11673" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11674" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7143" />
                    <RANKING order="2" place="2" resultid="7271" />
                    <RANKING order="3" place="3" resultid="6979" />
                    <RANKING order="4" place="4" resultid="7840" />
                    <RANKING order="5" place="5" resultid="7123" />
                    <RANKING order="6" place="6" resultid="9092" />
                    <RANKING order="7" place="7" resultid="6790" />
                    <RANKING order="8" place="8" resultid="7674" />
                    <RANKING order="9" place="-1" resultid="7817" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8626" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8627" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1504" daytime="11:45" gender="F" number="31" order="14" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11675" agemax="24" agemin="19" name="Pre-Masters">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6817" />
                    <RANKING order="2" place="2" resultid="6813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11676" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11677" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11678" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11679" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6838" />
                    <RANKING order="2" place="2" resultid="6971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11680" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11681" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11682" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11683" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11684" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11685" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11686" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11687" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11688" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11689" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11690" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11691" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11692" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11693" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11694" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7275" />
                    <RANKING order="2" place="2" resultid="6838" />
                    <RANKING order="3" place="3" resultid="6817" />
                    <RANKING order="4" place="4" resultid="6813" />
                    <RANKING order="5" place="5" resultid="7853" />
                    <RANKING order="6" place="6" resultid="6971" />
                    <RANKING order="7" place="7" resultid="7532" />
                    <RANKING order="8" place="-1" resultid="7218" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8628" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8629" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1522" daytime="11:55" gender="M" number="32" order="15" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11695" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11696" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11697" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11698" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7823" />
                    <RANKING order="2" place="2" resultid="6944" />
                    <RANKING order="3" place="3" resultid="7873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11699" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7268" />
                    <RANKING order="2" place="2" resultid="7198" />
                    <RANKING order="3" place="3" resultid="6937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11700" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6805" />
                    <RANKING order="2" place="2" resultid="9095" />
                    <RANKING order="3" place="-1" resultid="7244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11701" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11702" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7137" />
                    <RANKING order="2" place="2" resultid="6798" />
                    <RANKING order="3" place="-1" resultid="7234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11703" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11704" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11705" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="7249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11706" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11707" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11708" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11709" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11710" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11711" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11712" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11713" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11714" agemax="-1" agemin="-1" name="Klassierung nach Zeit">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7823" />
                    <RANKING order="2" place="2" resultid="6944" />
                    <RANKING order="3" place="3" resultid="7873" />
                    <RANKING order="4" place="4" resultid="7268" />
                    <RANKING order="5" place="5" resultid="6805" />
                    <RANKING order="6" place="6" resultid="7137" />
                    <RANKING order="7" place="7" resultid="7198" />
                    <RANKING order="8" place="8" resultid="7131" />
                    <RANKING order="9" place="9" resultid="6798" />
                    <RANKING order="10" place="10" resultid="6937" />
                    <RANKING order="11" place="11" resultid="7229" />
                    <RANKING order="12" place="12" resultid="9095" />
                    <RANKING order="13" place="-1" resultid="7244" />
                    <RANKING order="14" place="-1" resultid="7249" />
                    <RANKING order="15" place="-1" resultid="7234" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8630" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8631" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-27" daytime="12:10" name="Sonntag -- Staffeln" number="8">
          <EVENTS>
            <EVENT eventid="1540" daytime="12:10" gender="X" number="33" order="17" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="2000" />
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2001" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7433" />
                    <RANKING order="2" place="2" resultid="6883" />
                    <RANKING order="3" place="3" resultid="7291" />
                    <RANKING order="4" place="4" resultid="7011" />
                    <RANKING order="5" place="5" resultid="7438" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8633" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-27" name="Staffeln der Behinderten" number="9">
          <EVENTS>
            <EVENT eventid="7349" number="35" order="21" preveventid="-1" round="TIM">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7357" agemax="-1" agemin="-1" name="Behinderte (Klasse 20)" />
                <AGEGROUP agegroupid="7350" agemax="-1" agemin="-1" name="Behinderte (Klasse 34)" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="11716" number="34" order="20" preveventid="-1" round="TIM">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11718" agemax="-1" agemin="-1" name="Behinderte (Klasse 20)" />
                <AGEGROUP agegroupid="11719" agemax="-1" agemin="-1" name="Behinderte (Klasse 34)" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="WAED" name="Schwimmverein Wädenswil" nation="SUI" region="RZO">
          <CONTACT city="Wädenswil" name="Truttmann Otto" phone="044 780 75 06" street="Freiherrenstrasse 4" zip="8820" />
          <ATHLETES>
            <ATHLETE birthdate="1954-01-12" firstname="Ales" gender="M" lastname="Vrana" nation="SUI" license="19251" athleteid="6774">
              <RESULTS>
                <RESULT eventid="1414" points="712" swimtime="00:01:23.18" resultid="6777" lane="5" heatid="8614">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="702" swimtime="00:00:37.35" resultid="6775" lane="4" heatid="8547" />
                <RESULT eventid="1304" points="708" swimtime="00:03:04.84" resultid="6776" lane="1" heatid="8584">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:28.57" />
                    <SPLIT distance="150" swimtime="00:02:17.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SV 01" name="Mainzer SV 01" nation="GER">
          <CONTACT city="Mainz-Gonsenheim" country="DE" email="Guenter.Schmah@mainzersv01.de10" name="Schmah Günter" phone="06131-474854" state="RP" street="Max-Planck-Strasse 35c" zip="55124" />
          <ATHLETES>
            <ATHLETE birthdate="1938-01-01" firstname="Günter" gender="M" lastname="Schmah" nation="GER" license="12094" athleteid="6779">
              <RESULTS>
                <RESULT eventid="1342" points="485" swimtime="00:01:42.47" resultid="6784" lane="5" heatid="8600">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="787" swimtime="00:03:31.14" resultid="6783" lane="3" heatid="8583">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.23" />
                    <SPLIT distance="100" swimtime="00:01:43.69" />
                    <SPLIT distance="150" swimtime="00:02:38.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="504" swimtime="00:00:42.84" resultid="6782" lane="6" heatid="8559" />
                <RESULT eventid="1284" points="760" swimtime="00:00:41.88" resultid="6781" lane="5" heatid="8546" />
                <RESULT eventid="1414" points="806" swimtime="00:01:34.06" resultid="6785" lane="3" heatid="8613">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-01-01" firstname="Franz" gender="M" lastname="Schlömer" nation="GER" license="12095" athleteid="6780">
              <RESULTS>
                <RESULT eventid="1288" points="576" swimtime="00:01:36.04" resultid="6786" lane="4" heatid="8554">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="358" swimtime="00:01:46.33" resultid="6787" lane="1" heatid="8565">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="508" swimtime="00:03:38.71" resultid="6790" lane="3" heatid="8626">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.93" />
                    <SPLIT distance="100" swimtime="00:01:44.85" />
                    <SPLIT distance="150" swimtime="00:02:42.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="410" swimtime="00:01:49.60" resultid="6789" lane="2" heatid="8613">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="434" swimtime="00:00:46.58" resultid="6788" lane="3" heatid="8606" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCFG" name="SC Flipper Gossau" nation="SUI" region="ROS">
          <CONTACT city="Gossau" email="benedikt.rusch@helvetia.ch" fax="079 696 35 89" name="Rusch Benedikt" phone="058 280 43 65" street="Ilgenstrasse 7" zip="9200" />
          <ATHLETES>
            <ATHLETE birthdate="1954-01-01" firstname="Benedikt" gender="M" lastname="Rusch" nation="SUI" license="6282" athleteid="6792">
              <RESULTS>
                <RESULT eventid="1196" points="835" swimtime="00:10:38.32" resultid="6795" lane="1" heatid="8590">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                    <SPLIT distance="100" swimtime="00:01:15.15" />
                    <SPLIT distance="150" swimtime="00:01:55.54" />
                    <SPLIT distance="200" swimtime="00:02:36.28" />
                    <SPLIT distance="250" swimtime="00:03:17.45" />
                    <SPLIT distance="300" swimtime="00:03:58.73" />
                    <SPLIT distance="350" swimtime="00:04:39.86" />
                    <SPLIT distance="400" swimtime="00:05:20.98" />
                    <SPLIT distance="450" swimtime="00:06:01.07" />
                    <SPLIT distance="500" swimtime="00:06:41.11" />
                    <SPLIT distance="550" swimtime="00:07:20.66" />
                    <SPLIT distance="600" swimtime="00:08:00.47" />
                    <SPLIT distance="650" swimtime="00:08:40.16" />
                    <SPLIT distance="700" swimtime="00:09:20.09" />
                    <SPLIT distance="750" swimtime="00:10:00.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="647" swimtime="00:00:32.45" resultid="6794" lane="4" heatid="8559" />
                <RESULT comment="Schweizer Masters Rekord" eventid="1107" points="803" swimtime="00:02:21.75" resultid="6793" lane="2" heatid="8540">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:06.32" />
                    <SPLIT distance="150" swimtime="00:01:43.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="848" swimtime="00:05:02.42" resultid="6796" lane="3" heatid="8597">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:01:48.62" />
                    <SPLIT distance="200" swimtime="00:02:27.36" />
                    <SPLIT distance="250" swimtime="00:03:06.43" />
                    <SPLIT distance="300" swimtime="00:03:45.49" />
                    <SPLIT distance="350" swimtime="00:04:24.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1450" points="782" swimtime="00:01:03.69" resultid="6797" lane="5" heatid="8623">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1522" points="669" swimtime="00:02:56.88" resultid="6798" lane="2" heatid="8630">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:21.09" />
                    <SPLIT distance="150" swimtime="00:02:13.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SVE" name="Schwimmverein Emmen" nation="SUI" region="RZW">
          <ATHLETES>
            <ATHLETE birthdate="1962-10-12" firstname="Martin" gender="M" lastname="Grapentin" nation="SUI" license="25754" athleteid="6800">
              <RESULTS>
                <RESULT eventid="1522" points="698" swimtime="00:02:37.58" resultid="6805" lane="3" heatid="8630">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="100" swimtime="00:01:13.11" />
                    <SPLIT distance="150" swimtime="00:02:00.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="740" swimtime="00:00:27.11" resultid="6802" lane="2" heatid="8580" />
                <RESULT eventid="1292" points="871" swimtime="00:00:28.68" resultid="6801" lane="5" heatid="8561" />
                <RESULT eventid="1342" points="819" swimtime="00:01:05.56" resultid="6803" lane="1" heatid="8601">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UET" name="SC Delphin Uetendorf" nation="SUI">
          <CONTACT city="Wattenwil" name="Berger Marianne" phone="033 356 24 38" street="Stafelalpstr.12" zip="3665" />
          <ATHLETES>
            <ATHLETE birthdate="1985-11-22" firstname="Nadja" gender="F" lastname="Bigler" nation="SUI" license="10084" athleteid="6807">
              <RESULTS>
                <RESULT eventid="1282" points="587" swimtime="00:00:39.16" resultid="6808" lane="4" heatid="8544" />
                <RESULT eventid="1294" points="628" swimtime="00:01:18.21" resultid="6809" lane="4" heatid="8564">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="555" swimtime="00:01:25.84" resultid="6812" lane="3" heatid="8611">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="612" swimtime="00:02:58.94" resultid="6810" lane="3" heatid="8582">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:24.84" />
                    <SPLIT distance="150" swimtime="00:02:11.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="457" swimtime="00:05:29.10" resultid="6811" lane="2" heatid="8595">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:01:16.63" />
                    <SPLIT distance="150" swimtime="00:01:58.55" />
                    <SPLIT distance="200" swimtime="00:02:40.81" />
                    <SPLIT distance="250" swimtime="00:03:23.08" />
                    <SPLIT distance="300" swimtime="00:04:05.95" />
                    <SPLIT distance="350" swimtime="00:04:48.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="522" swimtime="00:02:52.54" resultid="6813" lane="2" heatid="8629">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:22.52" />
                    <SPLIT distance="150" swimtime="00:02:12.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-10-06" firstname="Andrea" gender="F" lastname="Brechbühl" nation="SUI" license="15382" athleteid="6814">
              <RESULTS>
                <RESULT eventid="1504" points="573" swimtime="00:02:47.18" resultid="6817" lane="5" heatid="8629">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:20.35" />
                    <SPLIT distance="150" swimtime="00:02:09.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="522" swimtime="00:05:14.82" resultid="6815" lane="6" heatid="8595">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="150" swimtime="00:01:52.13" />
                    <SPLIT distance="200" swimtime="00:02:31.94" />
                    <SPLIT distance="250" swimtime="00:03:12.22" />
                    <SPLIT distance="300" swimtime="00:03:52.67" />
                    <SPLIT distance="350" swimtime="00:04:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="536" swimtime="00:01:15.47" resultid="6816" lane="2" heatid="8599">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-28" firstname="Yves" gender="M" lastname="Marclay" nation="SUI" license="3121" athleteid="6818">
              <RESULTS>
                <RESULT eventid="1288" points="506" swimtime="00:01:11.11" resultid="6820" lane="2" heatid="8556">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="746" swimtime="00:00:32.47" resultid="6819" lane="1" heatid="8549" />
                <RESULT eventid="1300" points="593" swimtime="00:00:27.46" resultid="6822" lane="1" heatid="8581" />
                <RESULT eventid="1296" points="576" swimtime="00:01:10.01" resultid="6821" lane="6" heatid="8567">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCT" name="SC Thalwil" nation="SUI">
          <CONTACT city="Oberrieden" country="CH" email="heinzhaller@gmx.ch" name="Haller Heinz" street="Wiesengrundstr. 38" zip="8942" />
          <ATHLETES>
            <ATHLETE birthdate="1966-01-01" firstname="Robert" gender="M" lastname="Mundschin" nation="SUI" athleteid="6824">
              <RESULTS>
                <RESULT eventid="1292" points="534" swimtime="00:00:32.86" resultid="6898" lane="5" heatid="8560" />
                <RESULT eventid="1300" points="697" swimtime="00:00:27.54" resultid="6899" lane="3" heatid="8579" />
                <RESULT eventid="1450" points="642" swimtime="00:01:01.91" resultid="6902" lane="6" heatid="8623">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="569" swimtime="00:02:22.85" resultid="6897" lane="4" heatid="8540">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:01:10.53" />
                    <SPLIT distance="150" swimtime="00:01:47.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="523" swimtime="00:05:11.62" resultid="6900" lane="6" heatid="8598">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                    <SPLIT distance="150" swimtime="00:01:54.21" />
                    <SPLIT distance="200" swimtime="00:02:34.30" />
                    <SPLIT distance="250" swimtime="00:03:14.51" />
                    <SPLIT distance="300" swimtime="00:03:54.65" />
                    <SPLIT distance="350" swimtime="00:04:34.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="420" swimtime="00:00:37.39" resultid="6901" lane="1" heatid="8607" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Anja" gender="F" lastname="Gemperli" nation="SUI" athleteid="6887" />
            <ATHLETE birthdate="1959-01-01" firstname="Matthias" gender="M" lastname="Beusch" nation="SUI" athleteid="6888">
              <RESULTS>
                <RESULT eventid="1378" points="660" swimtime="00:00:35.16" resultid="6905" lane="6" heatid="8608" />
                <RESULT eventid="1292" points="671" swimtime="00:00:31.66" resultid="6904" lane="6" heatid="8561" />
                <RESULT eventid="1300" points="681" swimtime="00:00:28.83" resultid="6903" lane="3" heatid="8578" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Mauro" gender="M" lastname="Paulon" nation="SUI" athleteid="6889">
              <RESULTS>
                <RESULT eventid="1288" points="549" swimtime="00:01:11.79" resultid="6906" lane="2" heatid="8555">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="615" swimtime="00:00:27.22" resultid="6907" lane="4" heatid="8580" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Fritz" gender="M" lastname="Keller" nation="SUI" athleteid="6890">
              <RESULTS>
                <RESULT eventid="1450" points="285" swimtime="00:01:23.16" resultid="6911" lane="4" heatid="8621">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="366" swimtime="00:01:36.06" resultid="6910" lane="4" heatid="8613">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="352" swimtime="00:00:34.74" resultid="6909" lane="5" heatid="8576" />
                <RESULT eventid="1284" points="393" swimtime="00:00:41.93" resultid="6908" lane="6" heatid="8546" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Richard" gender="M" lastname="Niedermann" nation="SUI" athleteid="6891">
              <RESULTS>
                <RESULT eventid="1378" points="751" swimtime="00:00:33.68" resultid="6915" lane="3" heatid="8607" />
                <RESULT comment="Schweizer Masters Rekord" eventid="1288" points="750" swimtime="00:01:13.92" resultid="6912" lane="6" heatid="8556">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="712" swimtime="00:00:28.40" resultid="6914" lane="2" heatid="8579" />
                <RESULT comment="203 - Bewegen vor dem Startkommando" eventid="1296" status="DSQ" swimtime="00:01:14.33" resultid="6913" lane="5" heatid="8566">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Manuel" gender="M" lastname="Strickler" nation="SUI" athleteid="6892">
              <RESULTS>
                <RESULT eventid="1296" points="586" swimtime="00:01:13.74" resultid="6918" lane="2" heatid="8566">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="632" swimtime="00:01:18.25" resultid="6921" lane="3" heatid="8614">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="453" swimtime="00:01:19.07" resultid="6917" lane="5" heatid="8555">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="617" swimtime="00:00:34.64" resultid="6916" lane="1" heatid="8548" />
                <RESULT eventid="1378" points="464" swimtime="00:00:36.19" resultid="6920" lane="5" heatid="8607" />
                <RESULT eventid="1300" points="565" swimtime="00:00:29.53" resultid="6919" lane="4" heatid="8578" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Arthur" gender="M" lastname="Rösler" nation="SUI" athleteid="6893">
              <RESULTS>
                <RESULT eventid="1157" points="307" swimtime="00:07:04.14" resultid="6922" lane="3" heatid="8596">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:01:28.55" />
                    <SPLIT distance="150" swimtime="00:02:19.63" />
                    <SPLIT distance="200" swimtime="00:03:13.95" />
                    <SPLIT distance="250" swimtime="00:04:10.73" />
                    <SPLIT distance="300" swimtime="00:05:08.42" />
                    <SPLIT distance="350" swimtime="00:06:06.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Heinz" gender="M" lastname="Haller" nation="SUI" athleteid="6894">
              <RESULTS>
                <RESULT eventid="1284" points="654" swimtime="00:00:37.09" resultid="6923" lane="2" heatid="8547" />
                <RESULT comment="Schweizer Masters Rekord" eventid="1292" points="763" swimtime="00:00:30.34" resultid="6924" lane="4" heatid="8560" />
                <RESULT eventid="1300" points="649" swimtime="00:00:29.30" resultid="6925" lane="1" heatid="8578" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SV SS" name="Schwimmverein Sempachersee" nation="SUI">
          <CONTACT city="Willisau" country="CH" email="mcdiezi@bluemail.ch" name="Filli Martin" street="Höchhusmatt 19" zip="6030" />
          <ATHLETES>
            <ATHLETE birthdate="1939-01-01" firstname="Rene" gender="M" lastname="Diezi" nation="SUI" license="6098" athleteid="6826">
              <RESULTS>
                <RESULT eventid="1296" points="603" swimtime="00:01:31.31" resultid="6830" lane="2" heatid="8565">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Schweizer Masters Rekord" eventid="1288" points="667" swimtime="00:01:36.74" resultid="6829" lane="3" heatid="8554">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="674" swimtime="00:02:56.39" resultid="6828" lane="5" heatid="8539">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:24.08" />
                    <SPLIT distance="150" swimtime="00:02:10.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="633" swimtime="00:03:47.01" resultid="6831" lane="2" heatid="8583">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.51" />
                    <SPLIT distance="100" swimtime="00:01:48.36" />
                    <SPLIT distance="150" swimtime="00:02:48.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-01-01" firstname="Maya-Claire" gender="F" lastname="Diezi" nation="SUI" license="445" athleteid="6827">
              <RESULTS>
                <RESULT eventid="1177" points="344" swimtime="00:17:25.44" resultid="6834" lane="2" heatid="8587">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.48" />
                    <SPLIT distance="100" swimtime="00:01:59.53" />
                    <SPLIT distance="150" swimtime="00:03:04.88" />
                    <SPLIT distance="200" swimtime="00:04:09.85" />
                    <SPLIT distance="250" swimtime="00:05:18.11" />
                    <SPLIT distance="300" swimtime="00:06:23.83" />
                    <SPLIT distance="350" swimtime="00:07:32.27" />
                    <SPLIT distance="400" swimtime="00:08:38.15" />
                    <SPLIT distance="450" swimtime="00:09:45.84" />
                    <SPLIT distance="500" swimtime="00:10:51.19" />
                    <SPLIT distance="550" swimtime="00:11:58.39" />
                    <SPLIT distance="600" swimtime="00:13:04.80" />
                    <SPLIT distance="650" swimtime="00:14:09.56" />
                    <SPLIT distance="700" swimtime="00:15:16.43" />
                    <SPLIT distance="750" swimtime="00:16:20.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="477" swimtime="00:04:36.80" resultid="6833" lane="5" heatid="8582">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.37" />
                    <SPLIT distance="100" swimtime="00:02:13.10" />
                    <SPLIT distance="150" swimtime="00:03:23.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="360" swimtime="00:02:07.81" resultid="6832" lane="6" heatid="8563">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Simone" gender="F" lastname="Bürli" nation="SUI" athleteid="6926">
              <RESULTS>
                <RESULT eventid="1054" points="670" swimtime="00:02:23.76" resultid="6931" lane="5" heatid="8537">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:09.18" />
                    <SPLIT distance="150" swimtime="00:01:46.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1177" points="757" swimtime="00:10:14.67" resultid="6932" lane="4" heatid="8588">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                    <SPLIT distance="150" swimtime="00:01:50.78" />
                    <SPLIT distance="200" swimtime="00:02:29.29" />
                    <SPLIT distance="250" swimtime="00:03:08.06" />
                    <SPLIT distance="300" swimtime="00:03:46.82" />
                    <SPLIT distance="350" swimtime="00:04:25.33" />
                    <SPLIT distance="400" swimtime="00:05:03.83" />
                    <SPLIT distance="450" swimtime="00:05:42.31" />
                    <SPLIT distance="500" swimtime="00:06:20.71" />
                    <SPLIT distance="550" swimtime="00:06:59.54" />
                    <SPLIT distance="600" swimtime="00:07:38.34" />
                    <SPLIT distance="650" swimtime="00:08:17.22" />
                    <SPLIT distance="700" swimtime="00:08:56.48" />
                    <SPLIT distance="750" swimtime="00:09:35.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="662" swimtime="00:05:07.25" resultid="6933" lane="1" heatid="8595">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:53.93" />
                    <SPLIT distance="200" swimtime="00:02:32.88" />
                    <SPLIT distance="250" swimtime="00:03:11.73" />
                    <SPLIT distance="300" swimtime="00:03:50.58" />
                    <SPLIT distance="350" swimtime="00:04:29.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Martin" gender="M" lastname="Filli" nation="SUI" athleteid="6927">
              <RESULTS>
                <RESULT eventid="1296" points="417" swimtime="00:01:22.57" resultid="6934" lane="3" heatid="8565">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1522" points="387" swimtime="00:03:07.10" resultid="6937" lane="5" heatid="8630">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:34.08" />
                    <SPLIT distance="150" swimtime="00:02:26.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="451" swimtime="00:11:14.96" resultid="6935" lane="4" heatid="8589">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                    <SPLIT distance="100" swimtime="00:01:16.84" />
                    <SPLIT distance="150" swimtime="00:01:58.93" />
                    <SPLIT distance="200" swimtime="00:02:41.51" />
                    <SPLIT distance="250" swimtime="00:03:24.53" />
                    <SPLIT distance="300" swimtime="00:04:07.30" />
                    <SPLIT distance="350" swimtime="00:04:51.14" />
                    <SPLIT distance="400" swimtime="00:05:34.13" />
                    <SPLIT distance="450" swimtime="00:06:17.97" />
                    <SPLIT distance="500" swimtime="00:07:00.93" />
                    <SPLIT distance="550" swimtime="00:07:44.26" />
                    <SPLIT distance="600" swimtime="00:08:26.98" />
                    <SPLIT distance="650" swimtime="00:09:09.68" />
                    <SPLIT distance="700" swimtime="00:09:52.35" />
                    <SPLIT distance="750" swimtime="00:10:35.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1450" points="480" swimtime="00:01:08.19" resultid="6936" lane="5" heatid="8622">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="Brigitte" gender="F" lastname="Herzog" nation="SUI" athleteid="6928">
              <RESULTS>
                <RESULT eventid="1298" points="314" swimtime="00:00:39.98" resultid="6938" lane="3" heatid="8571" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Bruno" gender="M" lastname="Moll" nation="SUI" athleteid="6929">
              <RESULTS>
                <RESULT eventid="1300" points="728" swimtime="00:00:28.20" resultid="6939" lane="4" heatid="8576" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="Andreas" gender="M" lastname="Moll" nation="SUI" athleteid="6930">
              <RESULTS>
                <RESULT eventid="1300" points="283" swimtime="00:00:37.19" resultid="6940" lane="6" heatid="8576" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-16" firstname="Bertrand" gender="M" lastname="Grob" nation="SUI" athleteid="7878">
              <RESULTS>
                <RESULT eventid="1292" points="581" swimtime="00:00:30.12" resultid="7880" lane="3" heatid="8560" />
                <RESULT comment="203 - Bewegen vor dem Startkommando" eventid="1284" status="DSQ" swimtime="00:00:34.87" resultid="7879" lane="6" heatid="8548" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Heidi" gender="F" lastname="Arnold" nation="SUI" athleteid="8710" />
            <ATHLETE birthdate="1969-12-25" firstname="Andreas" gender="M" lastname="Murer" nation="SUI" athleteid="8711" />
            <ATHLETE firstname="Martin" gender="M" lastname="Grapentin" nation="SUI" athleteid="10220" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1175" swimtime="00:02:30.14" resultid="7437" lane="6" heatid="8585">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.18" />
                    <SPLIT distance="100" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:01:57.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6928" number="1" />
                    <RELAYPOSITION athleteid="7878" number="2" />
                    <RELAYPOSITION athleteid="6926" number="3" />
                    <RELAYPOSITION athleteid="6927" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1540" swimtime="00:02:12.28" resultid="7438" lane="1" heatid="8633">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6800" number="1" />
                    <RELAYPOSITION athleteid="6926" number="2" />
                    <RELAYPOSITION athleteid="8710" number="3" />
                    <RELAYPOSITION athleteid="6927" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1175" swimtime="00:03:11.09" resultid="7436" lane="1" heatid="8585">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.39" />
                    <SPLIT distance="100" swimtime="00:01:50.51" />
                    <SPLIT distance="150" swimtime="00:02:32.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6827" number="1" />
                    <RELAYPOSITION athleteid="8710" number="2" />
                    <RELAYPOSITION athleteid="6826" number="3" />
                    <RELAYPOSITION athleteid="8711" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="RFN" name="Red Fish Neuchatel" nation="SUI" region="RSR">
          <ATHLETES>
            <ATHLETE birthdate="1966-07-21" firstname="Claudia" gender="F" lastname="Lautenbacher" nation="SUI" athleteid="6836">
              <RESULTS>
                <RESULT eventid="1504" points="696" swimtime="00:02:46.71" resultid="6838" lane="4" heatid="8629">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:19.96" />
                    <SPLIT distance="150" swimtime="00:02:07.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="685" swimtime="00:01:25.21" resultid="6837" lane="4" heatid="8611">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-09-17" firstname="Philippe" gender="M" lastname="Allegrini" nation="SUI" license="2383" athleteid="7283">
              <RESULTS>
                <RESULT eventid="1196" points="906" swimtime="00:08:54.99" resultid="9741" lane="3" heatid="9736">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.55" />
                    <SPLIT distance="200" swimtime="00:02:08.97" />
                    <SPLIT distance="300" swimtime="00:03:16.24" />
                    <SPLIT distance="400" swimtime="00:04:23.82" />
                    <SPLIT distance="500" swimtime="00:05:30.99" />
                    <SPLIT distance="600" swimtime="00:06:38.18" />
                    <SPLIT distance="700" swimtime="00:07:45.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7347" points="1019" swimtime="00:16:54.68" resultid="7430" lane="4" heatid="8592">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="100" swimtime="00:01:02.55" />
                    <SPLIT distance="150" swimtime="00:01:35.50" />
                    <SPLIT distance="200" swimtime="00:02:08.97" />
                    <SPLIT distance="250" swimtime="00:02:42.61" />
                    <SPLIT distance="300" swimtime="00:03:16.24" />
                    <SPLIT distance="350" swimtime="00:03:49.86" />
                    <SPLIT distance="400" swimtime="00:04:23.82" />
                    <SPLIT distance="450" swimtime="00:04:57.36" />
                    <SPLIT distance="500" swimtime="00:05:30.99" />
                    <SPLIT distance="550" swimtime="00:06:04.66" />
                    <SPLIT distance="600" swimtime="00:06:38.18" />
                    <SPLIT distance="650" swimtime="00:07:11.90" />
                    <SPLIT distance="700" swimtime="00:07:45.95" />
                    <SPLIT distance="750" swimtime="00:08:20.40" />
                    <SPLIT distance="800" swimtime="00:08:54.99" />
                    <SPLIT distance="850" swimtime="00:09:29.19" />
                    <SPLIT distance="900" swimtime="00:10:03.53" />
                    <SPLIT distance="950" swimtime="00:10:38.06" />
                    <SPLIT distance="1000" swimtime="00:11:12.58" />
                    <SPLIT distance="1050" swimtime="00:11:47.02" />
                    <SPLIT distance="1100" swimtime="00:12:21.64" />
                    <SPLIT distance="1150" swimtime="00:12:56.41" />
                    <SPLIT distance="1200" swimtime="00:13:30.97" />
                    <SPLIT distance="1250" swimtime="00:14:04.98" />
                    <SPLIT distance="1300" swimtime="00:14:39.51" />
                    <SPLIT distance="1350" swimtime="00:15:13.98" />
                    <SPLIT distance="1400" swimtime="00:15:48.42" />
                    <SPLIT distance="1450" swimtime="00:16:22.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LN" name="Lausanne Natation" nation="SUI" region="RSR">
          <CONTACT city="Lausanne" email="cedric.cattaneo@gmail.com" fax="0216165160" name="Cattaneo Cédric" phone="0216165159" state="VD" street="Av. du Servan 32" zip="1006" />
          <ATHLETES>
            <ATHLETE birthdate="1984-07-04" firstname="Sébastien" gender="M" lastname="Boutinard Rouelle" nation="SUI" athleteid="6840">
              <RESULTS>
                <RESULT eventid="1378" points="447" swimtime="00:00:34.18" resultid="6842" lane="2" heatid="8606" />
                <RESULT eventid="1450" points="520" swimtime="00:01:02.86" resultid="6843" lane="6" heatid="8624">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="509" swimtime="00:00:28.47" resultid="6841" lane="1" heatid="8580" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-05-25" firstname="Rainer" gender="M" lastname="Buchholz" nation="GER" athleteid="6844">
              <RESULTS>
                <RESULT eventid="1300" points="770" swimtime="00:00:25.25" resultid="6846" lane="2" heatid="8581" />
                <RESULT eventid="1288" points="736" swimtime="00:01:05.11" resultid="6845" lane="4" heatid="8556">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1450" status="WDR" swimtime="00:00:00.00" resultid="6848" />
                <RESULT eventid="1378" status="WDR" swimtime="00:00:00.00" resultid="6847" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-26" firstname="Cédric" gender="M" lastname="Cattaneo" nation="SUI" athleteid="6849">
              <RESULTS>
                <RESULT eventid="1450" status="WDR" swimtime="00:00:00.00" resultid="6853" />
                <RESULT eventid="1414" status="WDR" swimtime="00:00:00.00" resultid="6852" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-05" firstname="Eavan" gender="F" lastname="Dorcey" nation="IRL" athleteid="6854" />
            <ATHLETE birthdate="1989-05-10" firstname="Agustin" gender="M" lastname="Gutierrez" nation="SUI" athleteid="6858">
              <RESULTS>
                <RESULT eventid="1450" points="510" swimtime="00:01:01.80" resultid="6862" lane="4" heatid="8623">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="516" swimtime="00:00:35.31" resultid="6859" lane="3" heatid="8547" />
                <RESULT eventid="1414" points="489" swimtime="00:01:18.87" resultid="6861" lane="2" heatid="8614">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="558" swimtime="00:00:27.10" resultid="6860" lane="4" heatid="8579" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-21" firstname="Osamu" gender="M" lastname="Moser" nation="SUI" athleteid="6863">
              <RESULTS>
                <RESULT eventid="1414" points="588" swimtime="00:01:15.42" resultid="6866" lane="1" heatid="8615">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="637" swimtime="00:01:07.30" resultid="6865" lane="5" heatid="8567">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="646" swimtime="00:00:32.71" resultid="6864" lane="5" heatid="8549" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-21" firstname="Nicole" gender="F" lastname="Solenthaler" nation="SUI" athleteid="6867">
              <RESULTS>
                <RESULT eventid="1360" points="398" swimtime="00:00:40.48" resultid="6871" lane="4" heatid="8604" />
                <RESULT eventid="1286" points="437" swimtime="00:01:24.41" resultid="6868" lane="4" heatid="8552">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="344" swimtime="00:01:19.62" resultid="6872" lane="4" heatid="8618">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="412" swimtime="00:01:30.03" resultid="6869" lane="1" heatid="8564">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="376" swimtime="00:00:35.46" resultid="6870" lane="1" heatid="8573" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-16" firstname="David" gender="M" lastname="Tron" nation="LUX" athleteid="6873">
              <RESULTS>
                <RESULT eventid="1378" points="531" swimtime="00:00:32.28" resultid="6876" lane="1" heatid="8608" />
                <RESULT eventid="1296" points="590" swimtime="00:01:09.03" resultid="6874" lane="1" heatid="8567">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1450" points="582" swimtime="00:01:00.56" resultid="6877" lane="2" heatid="8624">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="571" swimtime="00:00:27.40" resultid="6875" lane="6" heatid="8581" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-04-10" firstname="Moira" gender="F" lastname="Wacker" nation="SUI" athleteid="6878">
              <RESULTS>
                <RESULT eventid="1298" points="429" swimtime="00:00:33.94" resultid="6880" lane="4" heatid="8572" />
                <RESULT eventid="1396" points="426" swimtime="00:01:33.76" resultid="6881" lane="5" heatid="8611">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="480" swimtime="00:00:41.89" resultid="6879" lane="2" heatid="8544" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1175" swimtime="00:02:18.52" resultid="6882" lane="5" heatid="8585">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                    <SPLIT distance="100" swimtime="00:01:22.19" />
                    <SPLIT distance="150" swimtime="00:01:50.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6867" number="1" />
                    <RELAYPOSITION athleteid="6878" number="2" />
                    <RELAYPOSITION athleteid="6844" number="3" />
                    <RELAYPOSITION athleteid="6840" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1540" swimtime="00:02:02.02" resultid="6883" lane="2" heatid="8633">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6858" number="1" />
                    <RELAYPOSITION athleteid="6867" number="2" />
                    <RELAYPOSITION athleteid="6878" number="3" />
                    <RELAYPOSITION athleteid="6873" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AARE" name="Schwimmclub Aarefisch" nation="SUI">
          <CONTACT city="Aarau" email="samuel..nikles@bluewin.ch" street="Weihermattstr. 74/76" zip="5000" />
          <ATHLETES>
            <ATHLETE birthdate="1984-02-14" firstname="Samuel" gender="M" lastname="Niklès" nation="SUI" athleteid="6885">
              <RESULTS>
                <RESULT eventid="1300" points="269" swimtime="00:00:35.19" resultid="6886" lane="3" heatid="8575" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-04" firstname="Alfonso" gender="M" lastname="Die" nation="SUI" athleteid="8635">
              <RESULTS>
                <RESULT eventid="1300" points="395" swimtime="00:00:33.27" resultid="8656" lane="1" heatid="8574" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TMJPN" name="Tousuikai Masters" nation="JPN">
          <CONTACT city="Brugg" country="CH" email="Yohei.Sato@psi.ch" name="Yohei Sato" street="Sommerhaldenstrasse 1a" zip="5200" />
          <ATHLETES>
            <ATHLETE birthdate="1972-09-14" firstname="Yohei" gender="M" lastname="Sato" nation="JPN" license="13-110" athleteid="6942" externalid="720914-2">
              <RESULTS>
                <RESULT eventid="1522" points="637" swimtime="00:02:25.74" resultid="6944" lane="2" heatid="8631">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:08.94" />
                    <SPLIT distance="150" swimtime="00:01:50.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="572" swimtime="00:01:16.21" resultid="6943" lane="4" heatid="8614">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SVB" name="Schwimmverein beider Basel" nation="SUI" region="RZW">
          <CONTACT city="Therwil" email="mtolusso@hotmail.com" name="Tolusso Markus" phone="061 721 00 52" street="Teichstrasse 47" zip="4106" />
          <ATHLETES>
            <ATHLETE birthdate="1976-04-23" firstname="Peter" gender="M" lastname="Bezak" nation="SUI" license="279" athleteid="6946">
              <RESULTS>
                <RESULT eventid="1450" points="479" swimtime="00:01:04.69" resultid="6951" lane="2" heatid="8623">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="527" swimtime="00:00:31.26" resultid="6948" lane="1" heatid="8561" />
                <RESULT eventid="1157" points="475" swimtime="00:05:08.22" resultid="6950" lane="5" heatid="8598">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                    <SPLIT distance="150" swimtime="00:01:50.41" />
                    <SPLIT distance="200" swimtime="00:02:29.72" />
                    <SPLIT distance="250" swimtime="00:03:08.77" />
                    <SPLIT distance="300" swimtime="00:03:48.82" />
                    <SPLIT distance="350" swimtime="00:04:29.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="479" swimtime="00:00:29.48" resultid="6949" lane="2" heatid="8578" />
                <RESULT eventid="1284" points="487" swimtime="00:00:37.42" resultid="6947" lane="5" heatid="8547" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-09-17" firstname="Roger" gender="M" lastname="Birrer" nation="SUI" athleteid="6952">
              <RESULTS>
                <RESULT eventid="1378" points="824" swimtime="00:00:30.78" resultid="6957" lane="3" heatid="8608" />
                <RESULT eventid="1342" points="895" swimtime="00:01:03.64" resultid="6956" lane="4" heatid="8601">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-02" firstname="Stefan" gender="M" lastname="Brand" nation="SUI" license="8010" athleteid="6958">
              <RESULTS>
                <RESULT eventid="1292" points="872" swimtime="00:00:26.54" resultid="6959" lane="3" heatid="8561" />
                <RESULT eventid="1450" points="884" swimtime="00:00:52.69" resultid="6962" lane="3" heatid="8624">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="811" swimtime="00:00:59.56" resultid="6961" lane="3" heatid="8601">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="804" swimtime="00:00:24.45" resultid="6960" lane="4" heatid="8581" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Heidi" gender="F" lastname="Clark" nation="SUI" athleteid="6963">
              <RESULTS>
                <RESULT eventid="1298" points="470" swimtime="00:00:33.94" resultid="6965" lane="6" heatid="8573" />
                <RESULT eventid="1432" points="437" swimtime="00:01:15.70" resultid="7014" lane="1" heatid="8619">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="418" swimtime="00:05:55.72" resultid="7013" lane="4" heatid="8594">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:25.12" />
                    <SPLIT distance="150" swimtime="00:02:10.63" />
                    <SPLIT distance="200" swimtime="00:02:56.33" />
                    <SPLIT distance="250" swimtime="00:03:41.64" />
                    <SPLIT distance="300" swimtime="00:04:26.29" />
                    <SPLIT distance="350" swimtime="00:05:11.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1054" points="402" swimtime="00:02:46.43" resultid="6964" lane="4" heatid="8536">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="100" swimtime="00:01:20.51" />
                    <SPLIT distance="150" swimtime="00:02:04.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-03" firstname="Margarethe" gender="F" lastname="Denk" nation="GER" license="18490" athleteid="6966">
              <RESULTS>
                <RESULT eventid="1324" points="459" swimtime="00:01:25.13" resultid="6970" lane="5" heatid="8599">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1177" points="461" swimtime="00:12:12.32" resultid="6969" lane="5" heatid="8588">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:01:27.47" />
                    <SPLIT distance="150" swimtime="00:02:14.57" />
                    <SPLIT distance="200" swimtime="00:03:01.90" />
                    <SPLIT distance="250" swimtime="00:03:48.44" />
                    <SPLIT distance="300" swimtime="00:04:35.40" />
                    <SPLIT distance="350" swimtime="00:05:22.20" />
                    <SPLIT distance="400" swimtime="00:06:08.92" />
                    <SPLIT distance="450" swimtime="00:06:55.36" />
                    <SPLIT distance="500" swimtime="00:07:40.89" />
                    <SPLIT distance="550" swimtime="00:08:26.68" />
                    <SPLIT distance="600" swimtime="00:09:13.05" />
                    <SPLIT distance="650" swimtime="00:09:58.99" />
                    <SPLIT distance="700" swimtime="00:10:44.66" />
                    <SPLIT distance="750" swimtime="00:11:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="532" swimtime="00:01:24.36" resultid="6968" lane="5" heatid="8564">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="576" swimtime="00:00:35.63" resultid="6967" lane="4" heatid="8557" />
                <RESULT eventid="1504" points="500" swimtime="00:03:06.16" resultid="6971" lane="2" heatid="8628">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="100" swimtime="00:01:31.59" />
                    <SPLIT distance="150" swimtime="00:02:25.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-09-26" firstname="Kurt" gender="M" lastname="Frei" nation="SUI" license="4468" athleteid="6972">
              <RESULTS>
                <RESULT eventid="1486" points="856" swimtime="00:02:50.49" resultid="6979" lane="5" heatid="8627">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:24.30" />
                    <SPLIT distance="150" swimtime="00:02:08.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="788" swimtime="00:00:36.19" resultid="6978" lane="2" heatid="8607" />
                <RESULT eventid="1288" points="721" swimtime="00:01:22.06" resultid="6974" lane="1" heatid="8556">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="727" swimtime="00:05:28.13" resultid="6977" lane="2" heatid="8597">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:01:18.79" />
                    <SPLIT distance="150" swimtime="00:02:01.04" />
                    <SPLIT distance="200" swimtime="00:02:43.17" />
                    <SPLIT distance="250" swimtime="00:03:25.55" />
                    <SPLIT distance="300" swimtime="00:04:07.81" />
                    <SPLIT distance="350" swimtime="00:04:49.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="727" swimtime="00:11:14.92" resultid="6976" lane="3" heatid="8589">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:22.21" />
                    <SPLIT distance="150" swimtime="00:02:06.18" />
                    <SPLIT distance="200" swimtime="00:02:49.79" />
                    <SPLIT distance="250" swimtime="00:03:33.06" />
                    <SPLIT distance="300" swimtime="00:04:16.07" />
                    <SPLIT distance="350" swimtime="00:04:59.15" />
                    <SPLIT distance="400" swimtime="00:05:42.20" />
                    <SPLIT distance="450" swimtime="00:06:24.95" />
                    <SPLIT distance="500" swimtime="00:07:07.81" />
                    <SPLIT distance="550" swimtime="00:07:50.18" />
                    <SPLIT distance="600" swimtime="00:08:32.86" />
                    <SPLIT distance="650" swimtime="00:09:14.98" />
                    <SPLIT distance="700" swimtime="00:09:57.02" />
                    <SPLIT distance="750" swimtime="00:10:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="529" swimtime="00:00:33.74" resultid="6975" lane="5" heatid="8577" />
                <RESULT eventid="1107" points="611" swimtime="00:02:46.39" resultid="6973" lane="1" heatid="8540">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:20.04" />
                    <SPLIT distance="150" swimtime="00:02:03.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-10" firstname="Irene" gender="F" lastname="Nestor" nation="SUI" license="607" athleteid="6980">
              <RESULTS>
                <RESULT eventid="1286" points="773" swimtime="00:01:29.31" resultid="6982" lane="3" heatid="8551">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1054" points="618" swimtime="00:02:56.59" resultid="6981" lane="5" heatid="8536">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:01:27.27" />
                    <SPLIT distance="150" swimtime="00:02:12.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="495" swimtime="00:01:37.94" resultid="6983" lane="4" heatid="8563">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="863" swimtime="00:03:14.85" resultid="6987" lane="4" heatid="8625">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.97" />
                    <SPLIT distance="100" swimtime="00:01:35.85" />
                    <SPLIT distance="150" swimtime="00:02:25.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1177" points="740" swimtime="00:12:38.34" resultid="6984" lane="3" heatid="8587">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                    <SPLIT distance="150" swimtime="00:02:20.53" />
                    <SPLIT distance="200" swimtime="00:03:08.81" />
                    <SPLIT distance="250" swimtime="00:03:57.12" />
                    <SPLIT distance="300" swimtime="00:04:45.42" />
                    <SPLIT distance="350" swimtime="00:05:33.17" />
                    <SPLIT distance="400" swimtime="00:06:20.88" />
                    <SPLIT distance="450" swimtime="00:07:08.51" />
                    <SPLIT distance="500" swimtime="00:07:56.35" />
                    <SPLIT distance="550" swimtime="00:08:44.14" />
                    <SPLIT distance="600" swimtime="00:09:31.85" />
                    <SPLIT distance="650" swimtime="00:10:19.40" />
                    <SPLIT distance="700" swimtime="00:11:06.93" />
                    <SPLIT distance="750" swimtime="00:11:54.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="765" swimtime="00:06:04.60" resultid="6985" lane="1" heatid="8594">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                    <SPLIT distance="100" swimtime="00:01:29.99" />
                    <SPLIT distance="150" swimtime="00:02:17.04" />
                    <SPLIT distance="200" swimtime="00:03:03.53" />
                    <SPLIT distance="250" swimtime="00:03:49.63" />
                    <SPLIT distance="300" swimtime="00:04:35.47" />
                    <SPLIT distance="350" swimtime="00:05:21.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1360" points="595" swimtime="00:00:44.04" resultid="6986" lane="6" heatid="8604" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-12-14" firstname="Ferdy" gender="M" lastname="Polasek" nation="SUI" license="16664" athleteid="6988">
              <RESULTS>
                <RESULT eventid="1157" points="636" swimtime="00:05:12.05" resultid="6993" lane="1" heatid="8598">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:15.24" />
                    <SPLIT distance="150" swimtime="00:01:55.39" />
                    <SPLIT distance="200" swimtime="00:02:35.91" />
                    <SPLIT distance="250" swimtime="00:03:16.31" />
                    <SPLIT distance="300" swimtime="00:03:56.39" />
                    <SPLIT distance="350" swimtime="00:04:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="624" swimtime="00:02:25.43" resultid="6989" lane="3" heatid="8540">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:10.32" />
                    <SPLIT distance="150" swimtime="00:01:47.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="480" swimtime="00:00:41.11" resultid="6990" lane="3" heatid="8546" />
                <RESULT eventid="1196" points="627" swimtime="00:11:02.37" resultid="6992" lane="6" heatid="8590">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:01:16.45" />
                    <SPLIT distance="150" swimtime="00:01:57.70" />
                    <SPLIT distance="200" swimtime="00:02:39.39" />
                    <SPLIT distance="250" swimtime="00:03:21.03" />
                    <SPLIT distance="300" swimtime="00:04:02.65" />
                    <SPLIT distance="350" swimtime="00:04:44.77" />
                    <SPLIT distance="400" swimtime="00:05:27.14" />
                    <SPLIT distance="450" swimtime="00:06:09.69" />
                    <SPLIT distance="500" swimtime="00:06:51.93" />
                    <SPLIT distance="550" swimtime="00:07:34.40" />
                    <SPLIT distance="600" swimtime="00:08:16.42" />
                    <SPLIT distance="650" swimtime="00:08:59.17" />
                    <SPLIT distance="700" swimtime="00:09:41.04" />
                    <SPLIT distance="750" swimtime="00:10:23.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1450" points="628" swimtime="00:01:06.40" resultid="6994" lane="3" heatid="8622">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="599" swimtime="00:00:30.09" resultid="6991" lane="5" heatid="8578" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-05-30" firstname="Mireille" gender="F" lastname="Richter" nation="SUI" license="5930" athleteid="6995">
              <RESULTS>
                <RESULT eventid="1396" points="430" swimtime="00:01:54.47" resultid="6999" lane="2" heatid="8610">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.35" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Schweizer Masters Rekord" eventid="1054" points="680" swimtime="00:03:04.11" resultid="6996" lane="3" heatid="8535">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                    <SPLIT distance="100" swimtime="00:01:31.05" />
                    <SPLIT distance="150" swimtime="00:02:18.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="502" swimtime="00:03:55.18" resultid="6997" lane="4" heatid="8582">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.75" />
                    <SPLIT distance="100" swimtime="00:01:54.37" />
                    <SPLIT distance="150" swimtime="00:02:54.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1177" points="777" swimtime="00:13:04.04" resultid="9734" lane="5" heatid="8587">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.09" />
                    <SPLIT distance="200" swimtime="00:03:15.86" />
                    <SPLIT distance="300" swimtime="00:04:55.26" />
                    <SPLIT distance="400" swimtime="00:06:33.45" />
                    <SPLIT distance="500" swimtime="00:08:11.96" />
                    <SPLIT distance="600" swimtime="00:09:50.13" />
                    <SPLIT distance="700" swimtime="00:11:28.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7347" points="857" swimtime="00:24:21.65" resultid="8684" lane="3" heatid="8592">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.88" />
                    <SPLIT distance="100" swimtime="00:01:36.09" />
                    <SPLIT distance="150" swimtime="00:02:26.16" />
                    <SPLIT distance="200" swimtime="00:03:15.86" />
                    <SPLIT distance="250" swimtime="00:04:05.42" />
                    <SPLIT distance="300" swimtime="00:04:55.26" />
                    <SPLIT distance="350" swimtime="00:05:44.30" />
                    <SPLIT distance="400" swimtime="00:06:33.45" />
                    <SPLIT distance="450" swimtime="00:07:22.44" />
                    <SPLIT distance="500" swimtime="00:08:11.96" />
                    <SPLIT distance="550" swimtime="00:09:01.00" />
                    <SPLIT distance="600" swimtime="00:09:50.13" />
                    <SPLIT distance="650" swimtime="00:10:39.32" />
                    <SPLIT distance="700" swimtime="00:11:28.05" />
                    <SPLIT distance="750" swimtime="00:12:16.15" />
                    <SPLIT distance="800" swimtime="00:13:04.04" />
                    <SPLIT distance="850" swimtime="00:13:52.38" />
                    <SPLIT distance="900" swimtime="00:14:41.29" />
                    <SPLIT distance="950" swimtime="00:15:30.90" />
                    <SPLIT distance="1000" swimtime="00:16:20.43" />
                    <SPLIT distance="1050" swimtime="00:17:09.29" />
                    <SPLIT distance="1100" swimtime="00:17:58.32" />
                    <SPLIT distance="1150" swimtime="00:18:46.59" />
                    <SPLIT distance="1200" swimtime="00:19:34.86" />
                    <SPLIT distance="1250" swimtime="00:20:23.09" />
                    <SPLIT distance="1300" swimtime="00:21:11.70" />
                    <SPLIT distance="1350" swimtime="00:21:59.75" />
                    <SPLIT distance="1400" swimtime="00:22:47.63" />
                    <SPLIT distance="1450" swimtime="00:23:35.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-15" firstname="Regula" gender="F" lastname="Steiger" nation="SUI" license="514" athleteid="7000">
              <RESULTS>
                <RESULT eventid="1298" points="1109" swimtime="00:00:29.96" resultid="7002" lane="4" heatid="8573" />
                <RESULT eventid="1396" points="1022" swimtime="00:01:26.65" resultid="7003" lane="2" heatid="8611">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="934" swimtime="00:00:39.35" resultid="7001" lane="3" heatid="8544" />
                <RESULT eventid="1432" status="DNS" swimtime="00:00:00.00" resultid="7004" lane="5" heatid="8619" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-08-10" firstname="Markus" gender="M" lastname="Tolusso" nation="SUI" athleteid="7005">
              <RESULTS>
                <RESULT eventid="1288" points="462" swimtime="00:01:26.91" resultid="7006" lane="6" heatid="8555">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="507" swimtime="00:01:22.17" resultid="7008" lane="4" heatid="8565">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="557" swimtime="00:00:33.69" resultid="7007" lane="6" heatid="8560" />
                <RESULT eventid="1196" points="529" swimtime="00:11:40.76" resultid="7010" lane="2" heatid="8589">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:01:22.25" />
                    <SPLIT distance="150" swimtime="00:02:07.00" />
                    <SPLIT distance="200" swimtime="00:02:51.27" />
                    <SPLIT distance="250" swimtime="00:03:36.36" />
                    <SPLIT distance="300" swimtime="00:04:21.00" />
                    <SPLIT distance="350" swimtime="00:05:05.19" />
                    <SPLIT distance="400" swimtime="00:05:49.66" />
                    <SPLIT distance="450" swimtime="00:06:33.68" />
                    <SPLIT distance="500" swimtime="00:07:17.61" />
                    <SPLIT distance="550" swimtime="00:08:01.90" />
                    <SPLIT distance="600" swimtime="00:08:46.34" />
                    <SPLIT distance="650" swimtime="00:09:30.49" />
                    <SPLIT distance="700" swimtime="00:10:14.43" />
                    <SPLIT distance="750" swimtime="00:10:58.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="492" swimtime="00:00:32.12" resultid="7009" lane="3" heatid="8576" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1540" swimtime="00:02:05.72" resultid="7011" lane="4" heatid="8633">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6946" number="1" />
                    <RELAYPOSITION athleteid="6963" number="2" />
                    <RELAYPOSITION athleteid="6988" number="3" />
                    <RELAYPOSITION athleteid="6966" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1175" swimtime="00:02:18.20" resultid="7012" lane="4" heatid="8585">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:18.14" />
                    <SPLIT distance="150" swimtime="00:01:44.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6972" number="1" />
                    <RELAYPOSITION athleteid="7000" number="2" />
                    <RELAYPOSITION athleteid="6958" number="3" />
                    <RELAYPOSITION athleteid="6963" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SRM" name="SK Region Murten" nation="SUI" region="RSR">
          <CONTACT city="Murten" email="keiju@bluewin.ch" name="Herzig Heidi" street="Prehlstr. 35" zip="3280" />
          <ATHLETES>
            <ATHLETE birthdate="1966-04-17" firstname="Alexis" gender="M" lastname="Bögli" nation="SUI" license="12118" athleteid="7081">
              <RESULTS>
                <RESULT eventid="1284" points="702" swimtime="00:00:33.18" resultid="7082" lane="6" heatid="8549" />
                <RESULT eventid="1414" points="648" swimtime="00:01:17.63" resultid="7085" lane="5" heatid="8615">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="618" swimtime="00:04:54.88" resultid="7084" lane="2" heatid="8598">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                    <SPLIT distance="150" swimtime="00:01:45.62" />
                    <SPLIT distance="200" swimtime="00:02:23.18" />
                    <SPLIT distance="250" swimtime="00:03:01.03" />
                    <SPLIT distance="300" swimtime="00:03:39.67" />
                    <SPLIT distance="350" swimtime="00:04:18.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="612" swimtime="00:00:28.76" resultid="7083" lane="3" heatid="8580" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-07-30" firstname="Anita" gender="F" lastname="Zingg" nation="SUI" license="4769" athleteid="7086">
              <RESULTS>
                <RESULT eventid="1286" points="787" swimtime="00:01:19.20" resultid="7088" lane="3" heatid="8552">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1054" points="712" swimtime="00:02:34.45" resultid="7087" lane="1" heatid="8537">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:13.55" />
                    <SPLIT distance="150" swimtime="00:01:53.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" status="WDR" swimtime="00:00:00.00" resultid="7089" />
                <RESULT eventid="1432" status="WDR" swimtime="00:00:00.00" resultid="7090" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WITT" name="Schwimm-Club Wittenbach" nation="SUI" region="ROS">
          <CONTACT city="St.Gallen" email="gabschneider@gmx.net" name="Schneider Gabriel" street="Lukasstr.5" zip="9008" />
          <ATHLETES>
            <ATHLETE birthdate="1972-11-11" firstname="Matthias" gender="M" lastname="Baumberger" nation="SUI" license="23131" athleteid="7092">
              <RESULTS>
                <RESULT eventid="1450" status="WDR" swimtime="00:00:00.00" resultid="7096" />
                <RESULT eventid="1157" status="WDR" swimtime="00:00:00.00" resultid="7095" />
                <RESULT eventid="1300" status="WDR" swimtime="00:00:00.00" resultid="7094" />
                <RESULT eventid="1107" status="WDR" swimtime="00:00:00.00" resultid="7093" />
                <RESULT eventid="1292" status="WDR" swimtime="00:00:00.00" resultid="7097" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PLAN" name="CN Plan-les-Ouates" nation="SUI" region="RSR">
          <CONTACT city="Châtelaine" email="rascha54@yahoo.fr" name="Schallon Ralph" phone="022 796 79 83" street="av. de Crozet 12" street2="Directeur technique" zip="1219" />
          <ATHLETES>
            <ATHLETE birthdate="1953-06-12" firstname="Alexandre" gender="M" lastname="Barrena" nation="SUI" license="13184" athleteid="7099" />
            <ATHLETE birthdate="1965-07-13" firstname="Murielle" gender="F" lastname="Caillet Dayer" nation="SUI" license="1035" athleteid="7102">
              <RESULTS>
                <RESULT eventid="1286" points="413" swimtime="00:01:29.51" resultid="7103" lane="4" heatid="8551">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="458" swimtime="00:03:08.65" resultid="7107" lane="3" heatid="8625">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.04" />
                    <SPLIT distance="100" swimtime="00:01:32.34" />
                    <SPLIT distance="150" swimtime="00:02:21.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1360" points="403" swimtime="00:00:42.55" resultid="7106" lane="5" heatid="8604" />
                <RESULT eventid="1298" points="404" swimtime="00:00:36.79" resultid="7105" lane="6" heatid="8572" />
                <RESULT eventid="1294" points="419" swimtime="00:01:31.35" resultid="7104" lane="5" heatid="8563">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-12-23" firstname="Patricia" gender="F" lastname="Kamm" nation="SUI" license="24901" athleteid="7108">
              <RESULTS>
                <RESULT eventid="1177" points="624" swimtime="00:12:01.38" resultid="7110" lane="4" heatid="8587">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:23.16" />
                    <SPLIT distance="150" swimtime="00:02:08.44" />
                    <SPLIT distance="200" swimtime="00:02:54.55" />
                    <SPLIT distance="250" swimtime="00:03:40.86" />
                    <SPLIT distance="300" swimtime="00:04:27.29" />
                    <SPLIT distance="350" swimtime="00:05:12.31" />
                    <SPLIT distance="400" swimtime="00:05:58.18" />
                    <SPLIT distance="450" swimtime="00:06:44.59" />
                    <SPLIT distance="500" swimtime="00:07:30.52" />
                    <SPLIT distance="550" swimtime="00:08:15.87" />
                    <SPLIT distance="600" swimtime="00:09:01.89" />
                    <SPLIT distance="650" swimtime="00:09:47.53" />
                    <SPLIT distance="700" swimtime="00:10:33.04" />
                    <SPLIT distance="750" swimtime="00:11:18.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="593" swimtime="00:05:48.68" resultid="7111" lane="3" heatid="8593">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                    <SPLIT distance="100" swimtime="00:01:23.36" />
                    <SPLIT distance="150" swimtime="00:02:08.71" />
                    <SPLIT distance="200" swimtime="00:02:53.50" />
                    <SPLIT distance="250" swimtime="00:03:37.95" />
                    <SPLIT distance="300" swimtime="00:04:22.22" />
                    <SPLIT distance="350" swimtime="00:05:06.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="613" swimtime="00:01:14.78" resultid="7112" lane="5" heatid="8618">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="687" swimtime="00:01:22.87" resultid="7109" lane="2" heatid="8552">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-07-21" firstname="Nathalie" gender="F" lastname="Landenbergue" nation="SUI" license="1736" athleteid="7113">
              <RESULTS>
                <RESULT eventid="1298" points="441" swimtime="00:00:35.72" resultid="7116" lane="2" heatid="8572" />
                <RESULT eventid="1282" points="475" swimtime="00:00:43.60" resultid="7114" lane="5" heatid="8544" />
                <RESULT eventid="1432" points="478" swimtime="00:01:15.38" resultid="7118" lane="2" heatid="8618">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="558" swimtime="00:01:31.22" resultid="7117" lane="1" heatid="8611">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="444" swimtime="00:01:29.63" resultid="7115" lane="6" heatid="8564">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-08-15" firstname="Xavier" gender="M" lastname="Louis" nation="SUI" license="23189" athleteid="7119">
              <RESULTS>
                <RESULT eventid="1288" points="458" swimtime="00:01:18.75" resultid="7120" lane="4" heatid="8555">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="446" swimtime="00:02:57.34" resultid="7123" lane="1" heatid="8627">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                    <SPLIT distance="150" swimtime="00:02:11.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="493" swimtime="00:00:35.45" resultid="7122" lane="4" heatid="8607" />
                <RESULT eventid="1300" points="599" swimtime="00:00:28.96" resultid="7121" lane="6" heatid="8579" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-03" firstname="Antoine" gender="M" lastname="Mayerat" nation="SUI" license="26076" athleteid="7124">
              <RESULTS>
                <RESULT eventid="1522" points="727" swimtime="00:02:45.21" resultid="7131" lane="6" heatid="8631">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="100" swimtime="00:01:17.81" />
                    <SPLIT distance="150" swimtime="00:02:06.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="704" swimtime="00:01:10.98" resultid="7129" lane="6" heatid="8601">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="666" swimtime="00:10:49.12" resultid="7128" lane="4" heatid="8590">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                    <SPLIT distance="100" swimtime="00:01:11.30" />
                    <SPLIT distance="150" swimtime="00:01:50.03" />
                    <SPLIT distance="200" swimtime="00:02:29.03" />
                    <SPLIT distance="250" swimtime="00:03:08.65" />
                    <SPLIT distance="300" swimtime="00:03:48.88" />
                    <SPLIT distance="350" swimtime="00:04:29.58" />
                    <SPLIT distance="400" swimtime="00:05:10.30" />
                    <SPLIT distance="450" swimtime="00:05:52.10" />
                    <SPLIT distance="500" swimtime="00:06:34.04" />
                    <SPLIT distance="550" swimtime="00:07:16.67" />
                    <SPLIT distance="600" swimtime="00:07:59.30" />
                    <SPLIT distance="650" swimtime="00:08:42.15" />
                    <SPLIT distance="700" swimtime="00:09:25.42" />
                    <SPLIT distance="750" swimtime="00:10:08.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1450" points="703" swimtime="00:01:03.97" resultid="7130" lane="1" heatid="8624">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="675" swimtime="00:02:21.69" resultid="7125" lane="2" heatid="8541">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:08.12" />
                    <SPLIT distance="150" swimtime="00:01:45.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="696" swimtime="00:00:31.29" resultid="7126" lane="2" heatid="8560" />
                <RESULT eventid="1300" points="672" swimtime="00:00:28.96" resultid="7127" lane="1" heatid="8579" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-07-02" firstname="Ralph" gender="M" lastname="Schallon" nation="SUI" license="3101" athleteid="7132">
              <RESULTS>
                <RESULT comment="World Masters Rekord" eventid="1304" points="1157" swimtime="00:02:36.90" resultid="7135" lane="2" heatid="8584">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:01:55.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="1098" swimtime="00:01:12.01" resultid="7136" lane="6" heatid="8615">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Schweizer Masters Rekord" eventid="1284" points="1015" swimtime="00:00:33.04" resultid="7133" lane="2" heatid="8548" />
                <RESULT eventid="1522" points="915" swimtime="00:02:39.40" resultid="7137" lane="4" heatid="8630">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:21.28" />
                    <SPLIT distance="150" swimtime="00:02:02.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" status="WDR" swimtime="00:00:00.00" resultid="7134" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1540" swimtime="00:02:05.24" resultid="7291" lane="5" heatid="8633">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7119" number="1" />
                    <RELAYPOSITION athleteid="7108" number="2" />
                    <RELAYPOSITION athleteid="7113" number="3" />
                    <RELAYPOSITION athleteid="7124" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1175" swimtime="00:02:28.87" resultid="7292" lane="2" heatid="8585">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.43" />
                    <SPLIT distance="100" swimtime="00:01:19.44" />
                    <SPLIT distance="150" swimtime="00:01:53.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7102" number="1" />
                    <RELAYPOSITION athleteid="7132" number="2" />
                    <RELAYPOSITION athleteid="7119" number="3" />
                    <RELAYPOSITION athleteid="7113" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AVU" name="Avully Natation" nation="SUI" region="RSR">
          <CONTACT city="Sézegnin" name="Gaspoz Olivier" phone="022 756 20 94" street="33 rte du Creux-du-Loup" zip="1285" />
          <ATHLETES>
            <ATHLETE birthdate="1973-08-24" firstname="Laurent" gender="M" lastname="Thévenaz" nation="SUI" license="17578" athleteid="7139">
              <RESULTS>
                <RESULT eventid="1486" points="639" swimtime="00:02:27.65" resultid="7143" lane="2" heatid="8627">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                    <SPLIT distance="150" swimtime="00:01:49.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="620" swimtime="00:04:47.80" resultid="7142" lane="4" heatid="8598">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:06.09" />
                    <SPLIT distance="150" swimtime="00:01:41.43" />
                    <SPLIT distance="200" swimtime="00:02:17.86" />
                    <SPLIT distance="250" swimtime="00:02:54.82" />
                    <SPLIT distance="300" swimtime="00:03:32.11" />
                    <SPLIT distance="350" swimtime="00:04:10.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="572" swimtime="00:10:20.41" resultid="7141" lane="5" heatid="8590">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="100" swimtime="00:01:08.19" />
                    <SPLIT distance="150" swimtime="00:01:45.44" />
                    <SPLIT distance="200" swimtime="00:02:23.37" />
                    <SPLIT distance="250" swimtime="00:03:01.53" />
                    <SPLIT distance="300" swimtime="00:03:40.89" />
                    <SPLIT distance="350" swimtime="00:04:20.65" />
                    <SPLIT distance="400" swimtime="00:05:00.30" />
                    <SPLIT distance="450" swimtime="00:05:39.89" />
                    <SPLIT distance="500" swimtime="00:06:20.00" />
                    <SPLIT distance="550" swimtime="00:07:00.79" />
                    <SPLIT distance="600" swimtime="00:07:41.40" />
                    <SPLIT distance="650" swimtime="00:08:22.08" />
                    <SPLIT distance="700" swimtime="00:09:02.92" />
                    <SPLIT distance="750" swimtime="00:09:42.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="648" swimtime="00:02:14.20" resultid="7140" lane="5" heatid="8541">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                    <SPLIT distance="100" swimtime="00:01:03.23" />
                    <SPLIT distance="150" swimtime="00:01:38.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BREM" name="SC Region Bremgarten" nation="SUI" region="RZO">
          <CONTACT city="Bremgarten 2" email="info@scrb.ch" internet="www.scrb.ch" name="Andy Kempter" street2="Postfach 2123" zip="5620" />
          <ATHLETES>
            <ATHLETE birthdate="1957-07-30" firstname="Brigitte" gender="F" lastname="Christen" nation="SUI" license="22603" athleteid="7147">
              <RESULTS>
                <RESULT eventid="1298" points="236" swimtime="00:00:47.11" resultid="7149" lane="1" heatid="8571" />
                <RESULT eventid="1054" points="267" swimtime="00:03:42.27" resultid="7148" lane="4" heatid="8535">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.97" />
                    <SPLIT distance="100" swimtime="00:01:48.15" />
                    <SPLIT distance="150" swimtime="00:02:46.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Matthias" gender="M" lastname="Fehlmann" nation="SUI" athleteid="7150">
              <RESULTS>
                <RESULT eventid="1284" points="311" swimtime="00:00:41.74" resultid="7152" lane="6" heatid="8547" />
                <RESULT comment="203 - Bewegen vor dem Startkommando" eventid="1107" status="DSQ" swimtime="00:02:44.80" resultid="7151" lane="2" heatid="8538">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:18.00" />
                    <SPLIT distance="150" swimtime="00:02:00.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" status="WDR" swimtime="00:00:00.00" resultid="7153" lane="6" heatid="8577" />
                <RESULT eventid="1304" status="WDR" swimtime="00:00:00.00" resultid="7154" lane="6" heatid="8584" />
                <RESULT eventid="1414" status="WDR" swimtime="00:00:00.00" resultid="7155" />
                <RESULT eventid="1450" status="WDR" swimtime="00:00:00.00" resultid="7156" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-12-06" firstname="Andy" gender="M" lastname="Kempter" nation="SUI" athleteid="7157">
              <RESULTS>
                <RESULT eventid="1378" points="393" swimtime="00:00:41.78" resultid="7160" lane="4" heatid="8606" />
                <RESULT eventid="1450" points="369" swimtime="00:01:19.25" resultid="7161" lane="3" heatid="8621">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="308" swimtime="00:00:41.05" resultid="7158" lane="4" heatid="8558" />
                <RESULT eventid="1300" points="414" swimtime="00:00:34.03" resultid="7159" lane="2" heatid="8576" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-08-09" firstname="Melanie" gender="F" lastname="Lins" nation="SUI" athleteid="7162">
              <RESULTS>
                <RESULT eventid="1282" points="297" swimtime="00:00:54.03" resultid="7163" lane="4" heatid="8543" />
                <RESULT comment="203 - Bewegen vor dem Startkommando" eventid="1298" status="DSQ" swimtime="00:00:42.89" resultid="7164" lane="5" heatid="8571" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-02-21" firstname="Ruth" gender="F" lastname="Stierli" nation="SUI" license="22083" athleteid="7165">
              <RESULTS>
                <RESULT eventid="1302" points="325" swimtime="00:04:19.38" resultid="7167" lane="2" heatid="8582">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.59" />
                    <SPLIT distance="100" swimtime="00:02:01.91" />
                    <SPLIT distance="150" swimtime="00:03:11.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="379" swimtime="00:00:52.37" resultid="7166" lane="3" heatid="8543" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Paul" gender="M" lastname="Spadt" nation="SUI" athleteid="7872">
              <RESULTS>
                <RESULT eventid="1522" points="593" swimtime="00:02:29.23" resultid="7873" lane="5" heatid="8631">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="150" swimtime="00:01:55.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BUEL" name="Schwimmclub Bülach" nation="SUI" region="RZO">
          <CONTACT city="Windlach" email="tibi.kiss@bluewin.ch" name="Kiss Tibor" phone="01/862 6001" street="Raaterstr. 20" zip="8175" />
          <ATHLETES>
            <ATHLETE birthdate="1983-03-01" firstname="Andrea" gender="F" lastname="Bächli" nation="SUI" license="10378" athleteid="7169">
              <RESULTS>
                <RESULT eventid="1294" points="567" swimtime="00:01:19.20" resultid="7174" lane="2" heatid="8564">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1177" points="763" swimtime="00:10:07.99" resultid="7171" lane="3" heatid="8588">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:51.70" />
                    <SPLIT distance="200" swimtime="00:02:29.98" />
                    <SPLIT distance="250" swimtime="00:03:08.38" />
                    <SPLIT distance="300" swimtime="00:03:46.92" />
                    <SPLIT distance="350" swimtime="00:04:25.21" />
                    <SPLIT distance="400" swimtime="00:05:03.69" />
                    <SPLIT distance="450" swimtime="00:05:41.87" />
                    <SPLIT distance="500" swimtime="00:06:20.16" />
                    <SPLIT distance="550" swimtime="00:06:58.90" />
                    <SPLIT distance="600" swimtime="00:07:37.25" />
                    <SPLIT distance="650" swimtime="00:08:15.67" />
                    <SPLIT distance="700" swimtime="00:08:53.40" />
                    <SPLIT distance="750" swimtime="00:09:31.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="597" swimtime="00:01:08.21" resultid="7173" lane="4" heatid="8619">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1054" points="612" swimtime="00:02:24.75" resultid="7170" lane="4" heatid="8537">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                    <SPLIT distance="150" swimtime="00:01:48.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="691" swimtime="00:05:00.79" resultid="7172" lane="4" heatid="8595">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:12.29" />
                    <SPLIT distance="150" swimtime="00:01:50.01" />
                    <SPLIT distance="200" swimtime="00:02:28.09" />
                    <SPLIT distance="250" swimtime="00:03:06.03" />
                    <SPLIT distance="300" swimtime="00:03:44.48" />
                    <SPLIT distance="350" swimtime="00:04:22.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-10" firstname="Patrice" gender="M" lastname="Pellaton" nation="SUI" license="1722" athleteid="7175">
              <RESULTS>
                <RESULT eventid="1107" points="640" swimtime="00:02:08.39" resultid="7176" lane="4" heatid="8541">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                    <SPLIT distance="100" swimtime="00:00:59.79" />
                    <SPLIT distance="150" swimtime="00:01:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="880" swimtime="00:00:23.73" resultid="7178" lane="3" heatid="8581" />
                <RESULT eventid="1292" points="812" swimtime="00:00:27.18" resultid="7177" lane="2" heatid="8561" />
                <RESULT eventid="1450" points="831" swimtime="00:00:53.80" resultid="7180" lane="4" heatid="8624">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="605" swimtime="00:01:05.67" resultid="7179" lane="2" heatid="8601">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-10-14" firstname="Alfredo" gender="M" lastname="Prencipe" nation="GER" athleteid="7181">
              <RESULTS>
                <RESULT eventid="1450" points="592" swimtime="00:01:03.59" resultid="7182" lane="3" heatid="8623">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="HSV" name="HSV Medizin Magdeburg" nation="GER">
          <CONTACT city="Magdeburg" email="klesinski@email.de" name="Gerald Schmidt" street="Hannoversche Str. 7d" zip="39110" />
          <ATHLETES>
            <ATHLETE birthdate="1976-09-22" firstname="René" gender="M" lastname="Klesinski" nation="GER" license="074167" athleteid="7184">
              <RESULTS>
                <RESULT eventid="1107" points="504" swimtime="00:02:20.31" resultid="7185" lane="1" heatid="8541">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:07.93" />
                    <SPLIT distance="150" swimtime="00:01:44.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="492" swimtime="00:00:31.99" resultid="7187" lane="2" heatid="8559" />
                <RESULT eventid="1288" points="402" swimtime="00:01:16.73" resultid="7186" lane="3" heatid="8555">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="431" swimtime="00:00:30.53" resultid="7188" lane="5" heatid="8579" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AMT" name="Aquatic Masters Team" nation="SUI">
          <CONTACT city="Bollingen" email="cristian58@bluewin.ch" name="Cristian Rentsch" street="Dorfstrasse 55" zip="8715" />
          <ATHLETES>
            <ATHLETE birthdate="1969-01-01" firstname="Basil" gender="M" lastname="Düby" nation="SUI" athleteid="7190">
              <RESULTS>
                <RESULT eventid="1342" points="586" swimtime="00:01:10.09" resultid="7196" lane="5" heatid="8601">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1522" points="611" swimtime="00:02:40.67" resultid="7198" lane="1" heatid="8631">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="100" swimtime="00:01:16.13" />
                    <SPLIT distance="150" swimtime="00:02:03.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1450" points="588" swimtime="00:01:03.74" resultid="7197" lane="1" heatid="8623">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Toni" gender="M" lastname="Pavicic-Donkic" nation="SUI" license="10982" athleteid="7191">
              <RESULTS>
                <RESULT eventid="1107" points="892" swimtime="00:02:02.95" resultid="7199" lane="3" heatid="8541">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                    <SPLIT distance="100" swimtime="00:00:59.19" />
                    <SPLIT distance="150" swimtime="00:01:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="916" swimtime="00:04:18.59" resultid="7267" lane="3" heatid="8598">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="100" swimtime="00:01:03.49" />
                    <SPLIT distance="150" swimtime="00:01:36.34" />
                    <SPLIT distance="200" swimtime="00:02:09.21" />
                    <SPLIT distance="250" swimtime="00:02:41.82" />
                    <SPLIT distance="300" swimtime="00:03:14.49" />
                    <SPLIT distance="350" swimtime="00:03:46.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1522" points="752" swimtime="00:02:29.93" resultid="7268" lane="4" heatid="8631">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="150" swimtime="00:01:54.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" status="DNS" swimtime="00:00:00.00" resultid="7266" lane="3" heatid="8590" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Christian" gender="M" lastname="Rentsch" nation="SUI" license="843" athleteid="7192">
              <RESULTS>
                <RESULT eventid="1304" points="856" swimtime="00:02:42.13" resultid="7270" lane="4" heatid="8584">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:18.17" />
                    <SPLIT distance="150" swimtime="00:02:00.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="846" swimtime="00:02:29.00" resultid="7271" lane="3" heatid="8627">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                    <SPLIT distance="100" swimtime="00:01:12.07" />
                    <SPLIT distance="150" swimtime="00:01:50.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="758" swimtime="00:00:33.69" resultid="7269" lane="4" heatid="8548" />
                <RESULT eventid="1157" status="DNS" swimtime="00:00:00.00" resultid="7662" lane="4" heatid="8597" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Sonja" gender="F" lastname="Gwerder" nation="SUI" license="13520" athleteid="7193">
              <RESULTS>
                <RESULT eventid="1504" points="684" swimtime="00:02:41.29" resultid="7275" lane="3" heatid="8629">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:16.76" />
                    <SPLIT distance="150" swimtime="00:02:03.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="830" swimtime="00:01:12.02" resultid="7272" lane="3" heatid="8564">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="732" swimtime="00:01:11.62" resultid="7273" lane="4" heatid="8599">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1360" points="854" swimtime="00:00:32.99" resultid="7274" lane="3" heatid="8604" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Alicia" gender="F" lastname="Irvin" nation="SUI" license="13815" athleteid="7194">
              <RESULTS>
                <RESULT eventid="1298" points="762" swimtime="00:00:29.34" resultid="7277" lane="3" heatid="8573" />
                <RESULT eventid="1054" points="423" swimtime="00:02:47.52" resultid="7276" lane="2" heatid="8536">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:21.13" />
                    <SPLIT distance="150" swimtime="00:02:04.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Evgenia" gender="F" lastname="Bedenig" nation="SUI" athleteid="7195">
              <RESULTS>
                <RESULT eventid="1290" points="452" swimtime="00:00:37.56" resultid="7279" lane="3" heatid="8557" />
                <RESULT eventid="1324" points="447" swimtime="00:01:23.66" resultid="7281" lane="3" heatid="8599">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="495" swimtime="00:01:13.38" resultid="7282" lane="3" heatid="8619">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1054" points="543" swimtime="00:02:33.52" resultid="7278" lane="3" heatid="8537">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:11.74" />
                    <SPLIT distance="150" swimtime="00:01:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="582" swimtime="00:05:20.97" resultid="7280" lane="3" heatid="8595">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:01:15.55" />
                    <SPLIT distance="150" swimtime="00:01:55.92" />
                    <SPLIT distance="200" swimtime="00:02:36.20" />
                    <SPLIT distance="250" swimtime="00:03:16.47" />
                    <SPLIT distance="300" swimtime="00:03:56.53" />
                    <SPLIT distance="350" swimtime="00:04:38.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <RESULTS>
                <RESULT eventid="1175" swimtime="00:02:05.44" resultid="7434" lane="3" heatid="8585">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                    <SPLIT distance="150" swimtime="00:01:36.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7192" number="1" />
                    <RELAYPOSITION athleteid="7191" number="2" />
                    <RELAYPOSITION athleteid="7193" number="3" />
                    <RELAYPOSITION athleteid="7194" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1540" swimtime="00:01:59.84" resultid="7433" lane="3" heatid="8633">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7190" number="1" />
                    <RELAYPOSITION athleteid="7191" number="2" />
                    <RELAYPOSITION athleteid="7193" number="3" />
                    <RELAYPOSITION athleteid="7195" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TSV" name="TSV 1862 Erding" nation="GER">
          <CONTACT email="delphine.erding@t-online.de" name="Petra Teichert" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Hans Georg" gender="M" lastname="Fiedeldeij" nation="GER" license="154290" athleteid="7201">
              <RESULTS>
                <RESULT eventid="1196" points="487" swimtime="00:10:57.90" resultid="7262" lane="2" heatid="8590">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:55.31" />
                    <SPLIT distance="200" swimtime="00:02:36.01" />
                    <SPLIT distance="250" swimtime="00:03:17.29" />
                    <SPLIT distance="300" swimtime="00:03:58.71" />
                    <SPLIT distance="350" swimtime="00:04:40.30" />
                    <SPLIT distance="400" swimtime="00:05:22.08" />
                    <SPLIT distance="450" swimtime="00:06:03.40" />
                    <SPLIT distance="500" swimtime="00:06:45.06" />
                    <SPLIT distance="550" swimtime="00:07:26.87" />
                    <SPLIT distance="600" swimtime="00:08:09.04" />
                    <SPLIT distance="650" swimtime="00:08:51.57" />
                    <SPLIT distance="700" swimtime="00:09:34.25" />
                    <SPLIT distance="750" swimtime="00:10:16.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="639" swimtime="00:00:28.34" resultid="7261" lane="5" heatid="8580" />
                <RESULT eventid="1107" points="528" swimtime="00:02:26.39" resultid="7260" lane="6" heatid="8541">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="100" swimtime="00:01:06.11" />
                    <SPLIT distance="150" swimtime="00:01:45.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCW" name="SC Winterthur" nation="SUI">
          <CONTACT email="mueller.peter@bluewin.ch" name="Peter Müller" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Markus" gender="M" lastname="Enz" nation="SUI" license="715" athleteid="7203">
              <RESULTS>
                <RESULT eventid="1296" points="566" swimtime="00:01:19.18" resultid="7255" lane="1" heatid="8566">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="594" swimtime="00:02:27.86" resultid="7252" lane="6" heatid="8540">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                    <SPLIT distance="100" swimtime="00:01:10.32" />
                    <SPLIT distance="150" swimtime="00:01:49.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="420" swimtime="00:00:37.00" resultid="7254" lane="5" heatid="8559" />
                <RESULT eventid="1300" points="560" swimtime="00:00:30.77" resultid="7256" lane="6" heatid="8578" />
                <RESULT comment="303 - Nicht mit beiden Händen gleich-zeitig angeschlagen (Wende  ...)" eventid="1284" status="DSQ" swimtime="00:00:38.12" resultid="7253" lane="1" heatid="8547" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Marcel" gender="M" lastname="Schwarz" nation="SUI" license="8657" athleteid="7204">
              <RESULTS>
                <RESULT eventid="1284" points="668" swimtime="00:00:32.36" resultid="7257" lane="3" heatid="8548" />
                <RESULT eventid="1300" points="585" swimtime="00:00:27.19" resultid="7259" lane="6" heatid="8580" />
                <RESULT comment="203 - Bewegen vor dem Startkommando" eventid="1296" status="DSQ" swimtime="00:01:06.56" resultid="7258" lane="2" heatid="8567">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNN" name="Cercle des Nageurs de Nyon" nation="SUI">
          <CONTACT city="Trelex" email="phil55@bluewin.ch" name="Mayer Philippe" phone="079 341 88 12" street="Chemin du treizou 7" zip="1270" />
          <ATHLETES>
            <ATHLETE birthdate="1955-01-01" firstname="Philippe" gender="M" lastname="Mayer" nation="SUI" license="4861" athleteid="7206">
              <RESULTS>
                <RESULT eventid="7347" points="579" swimtime="00:21:54.27" resultid="7431" lane="2" heatid="8592">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:01:59.54" />
                    <SPLIT distance="200" swimtime="00:02:40.36" />
                    <SPLIT distance="250" swimtime="00:03:22.77" />
                    <SPLIT distance="300" swimtime="00:04:05.32" />
                    <SPLIT distance="350" swimtime="00:04:48.20" />
                    <SPLIT distance="400" swimtime="00:05:31.66" />
                    <SPLIT distance="450" swimtime="00:06:16.27" />
                    <SPLIT distance="500" swimtime="00:07:00.42" />
                    <SPLIT distance="550" swimtime="00:07:44.21" />
                    <SPLIT distance="600" swimtime="00:08:28.28" />
                    <SPLIT distance="650" swimtime="00:09:12.36" />
                    <SPLIT distance="700" swimtime="00:09:55.73" />
                    <SPLIT distance="750" swimtime="00:10:38.62" />
                    <SPLIT distance="800" swimtime="00:11:22.01" />
                    <SPLIT distance="850" swimtime="00:12:15.09" />
                    <SPLIT distance="900" swimtime="00:13:02.07" />
                    <SPLIT distance="950" swimtime="00:13:48.29" />
                    <SPLIT distance="1000" swimtime="00:14:34.09" />
                    <SPLIT distance="1050" swimtime="00:15:19.14" />
                    <SPLIT distance="1100" swimtime="00:16:03.97" />
                    <SPLIT distance="1150" swimtime="00:16:48.67" />
                    <SPLIT distance="1200" swimtime="00:17:33.97" />
                    <SPLIT distance="1250" swimtime="00:18:18.57" />
                    <SPLIT distance="1300" swimtime="00:19:03.34" />
                    <SPLIT distance="1350" swimtime="00:19:47.33" />
                    <SPLIT distance="1400" swimtime="00:20:31.11" />
                    <SPLIT distance="1450" swimtime="00:21:14.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="574" swimtime="00:11:22.01" resultid="9740" lane="2" heatid="9736">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="200" swimtime="00:02:40.36" />
                    <SPLIT distance="300" swimtime="00:04:05.32" />
                    <SPLIT distance="400" swimtime="00:05:31.66" />
                    <SPLIT distance="500" swimtime="00:07:00.42" />
                    <SPLIT distance="600" swimtime="00:08:28.28" />
                    <SPLIT distance="700" swimtime="00:09:55.73" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="203 - Bewegen vor dem Startkommando" eventid="1304" status="DSQ" swimtime="00:02:45.86" resultid="7250" lane="5" heatid="8584">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:18.74" />
                    <SPLIT distance="150" swimtime="00:02:01.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOPR" name="Sport Figielski WOPR" nation="POL">
          <CONTACT country="PL" email="sport-figielski@02.pl" name="Grzegorz Figielski" />
          <ATHLETES>
            <ATHLETE birthdate="1958-01-01" firstname="Aleksandra" gender="F" lastname="Niespodziana" nation="POL" athleteid="7208">
              <RESULTS>
                <RESULT eventid="1504" status="WDR" swimtime="00:00:00.00" resultid="7218" />
                <RESULT eventid="1054" status="WDR" swimtime="00:00:00.00" resultid="7214" />
                <RESULT eventid="1290" status="WDR" swimtime="00:00:00.00" resultid="7215" />
                <RESULT eventid="1072" status="WDR" swimtime="00:00:00.00" resultid="7216" />
                <RESULT eventid="1324" status="WDR" swimtime="00:00:00.00" resultid="7217" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Grzegorz" gender="M" lastname="Figielski" nation="POL" athleteid="7210">
              <RESULTS>
                <RESULT eventid="1107" status="WDR" swimtime="00:00:00.00" resultid="7230" />
                <RESULT eventid="1196" status="WDR" swimtime="00:00:00.00" resultid="7231" />
                <RESULT eventid="1157" status="WDR" swimtime="00:00:00.00" resultid="7232" />
                <RESULT eventid="1342" status="WDR" swimtime="00:00:00.00" resultid="7233" />
                <RESULT eventid="1522" status="WDR" swimtime="00:00:00.00" resultid="7234" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="7211">
              <RESULTS>
                <RESULT eventid="1342" points="414" swimtime="00:01:24.73" resultid="7239" lane="4" heatid="8600">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7347" points="427" swimtime="00:24:14.40" resultid="8634" lane="5" heatid="8592">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:01:27.04" />
                    <SPLIT distance="150" swimtime="00:02:13.20" />
                    <SPLIT distance="200" swimtime="00:03:00.29" />
                    <SPLIT distance="250" swimtime="00:03:48.05" />
                    <SPLIT distance="300" swimtime="00:04:35.72" />
                    <SPLIT distance="350" swimtime="00:05:23.74" />
                    <SPLIT distance="400" swimtime="00:06:11.49" />
                    <SPLIT distance="450" swimtime="00:06:59.70" />
                    <SPLIT distance="500" swimtime="00:07:46.93" />
                    <SPLIT distance="550" swimtime="00:08:35.72" />
                    <SPLIT distance="600" swimtime="00:09:23.72" />
                    <SPLIT distance="650" swimtime="00:10:12.42" />
                    <SPLIT distance="700" swimtime="00:11:01.46" />
                    <SPLIT distance="750" swimtime="00:11:50.19" />
                    <SPLIT distance="800" swimtime="00:12:38.97" />
                    <SPLIT distance="850" swimtime="00:13:27.41" />
                    <SPLIT distance="900" swimtime="00:14:16.16" />
                    <SPLIT distance="950" swimtime="00:15:05.30" />
                    <SPLIT distance="1000" swimtime="00:15:53.69" />
                    <SPLIT distance="1050" swimtime="00:16:41.37" />
                    <SPLIT distance="1100" swimtime="00:17:29.58" />
                    <SPLIT distance="1150" swimtime="00:18:17.32" />
                    <SPLIT distance="1200" swimtime="00:19:05.80" />
                    <SPLIT distance="1250" swimtime="00:19:54.41" />
                    <SPLIT distance="1300" swimtime="00:20:42.39" />
                    <SPLIT distance="1350" swimtime="00:21:30.23" />
                    <SPLIT distance="1400" swimtime="00:22:18.02" />
                    <SPLIT distance="1450" swimtime="00:23:05.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="439" swimtime="00:02:43.46" resultid="7235" lane="3" heatid="8539">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:01:19.24" />
                    <SPLIT distance="150" swimtime="00:02:02.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="417" swimtime="00:12:38.97" resultid="9743" lane="4" heatid="9736">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.04" />
                    <SPLIT distance="200" swimtime="00:03:00.29" />
                    <SPLIT distance="300" swimtime="00:04:35.72" />
                    <SPLIT distance="400" swimtime="00:06:11.49" />
                    <SPLIT distance="500" swimtime="00:07:46.93" />
                    <SPLIT distance="600" swimtime="00:09:23.72" />
                    <SPLIT distance="700" swimtime="00:11:01.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="390" swimtime="00:00:37.93" resultid="8532" lane="1" heatid="8559" />
                <RESULT eventid="1300" points="451" swimtime="00:00:33.06" resultid="8531" lane="2" heatid="8577" />
                <RESULT eventid="1450" status="DNS" swimtime="00:00:00.00" resultid="8533" lane="2" heatid="8622" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Jacek" gender="M" lastname="Adamski" nation="POL" athleteid="7212">
              <RESULTS>
                <RESULT eventid="1522" status="WDR" swimtime="00:00:00.00" resultid="7244" />
                <RESULT eventid="1414" status="WDR" swimtime="00:00:00.00" resultid="7243" />
                <RESULT eventid="1296" status="WDR" swimtime="00:00:00.00" resultid="7241" />
                <RESULT eventid="1304" status="WDR" swimtime="00:00:00.00" resultid="7242" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-01-01" firstname="Zygmunt" gender="M" lastname="Lewandowski" nation="POL" athleteid="7213">
              <RESULTS>
                <RESULT eventid="1196" status="WDR" swimtime="00:00:00.00" resultid="7246" />
                <RESULT eventid="1522" status="WDR" swimtime="00:00:00.00" resultid="7249" />
                <RESULT eventid="1342" status="WDR" swimtime="00:00:00.00" resultid="7248" />
                <RESULT eventid="1296" status="WDR" swimtime="00:00:00.00" resultid="7245" />
                <RESULT eventid="1157" status="WDR" swimtime="00:00:00.00" resultid="7247" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SVZ" name="Schwimmverein Zürileu" nation="SUI" region="RZO">
          <CONTACT city="Urdorf" email="billabongs@gmx.net" internet="www.svzuerileu.ch" name="Axel Mathis-Pairo" phone="+41 79 404 31 35" state="SUI" street="Untermatt 5" zip="8902" />
          <ATHLETES>
            <ATHLETE birthdate="1959-06-16" firstname="Heike" gender="F" lastname="Lischke" nation="GER" license="25770" athleteid="7288">
              <RESULTS>
                <RESULT eventid="1396" points="662" swimtime="00:01:35.60" resultid="7289" lane="6" heatid="8611">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="415" swimtime="00:01:27.19" resultid="7290" lane="3" heatid="8617">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SKL" name="Schwimmklub Luzern" nation="SUI">
          <CONTACT city="Horw" name="Krejci Josef" phone="041 340 33 42" street="Stegenstrasse 29" zip="6048" />
          <ATHLETES>
            <ATHLETE birthdate="1936-11-17" firstname="Olga" gender="F" lastname="Krejci" nation="SUI" license="2600" athleteid="7294">
              <RESULTS>
                <RESULT eventid="1298" points="890" swimtime="00:00:39.16" resultid="7301" lane="4" heatid="8571" />
                <RESULT eventid="1282" points="635" swimtime="00:00:51.80" resultid="7300" lane="2" heatid="8543" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1933-05-18" firstname="Josef" gender="M" lastname="Krejci" nation="SUI" license="5618" athleteid="7295">
              <RESULTS>
                <RESULT comment="Schweizer Masters Rekord" eventid="1107" points="939" swimtime="00:02:53.27" resultid="7296" lane="3" heatid="8538">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:21.74" />
                    <SPLIT distance="150" swimtime="00:02:07.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="1113" swimtime="00:12:36.49" resultid="7297" lane="1" heatid="8589">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                    <SPLIT distance="100" swimtime="00:01:27.22" />
                    <SPLIT distance="150" swimtime="00:02:14.90" />
                    <SPLIT distance="200" swimtime="00:03:02.44" />
                    <SPLIT distance="250" swimtime="00:03:50.62" />
                    <SPLIT distance="300" swimtime="00:04:38.95" />
                    <SPLIT distance="350" swimtime="00:05:27.47" />
                    <SPLIT distance="400" swimtime="00:06:14.67" />
                    <SPLIT distance="450" swimtime="00:07:03.43" />
                    <SPLIT distance="500" swimtime="00:07:51.52" />
                    <SPLIT distance="550" swimtime="00:08:39.30" />
                    <SPLIT distance="600" swimtime="00:09:27.47" />
                    <SPLIT distance="650" swimtime="00:10:14.76" />
                    <SPLIT distance="700" swimtime="00:11:03.21" />
                    <SPLIT distance="750" swimtime="00:11:51.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DUCKS" name="Duck&apos;s Creek" nation="RUS">
          <CONTACT email="info@dcsport.ru" name="Vera Tarasova" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Vladislav" gender="M" lastname="Bragin" nation="RUS" athleteid="7333">
              <RESULTS>
                <RESULT eventid="1296" points="970" swimtime="00:00:58.99" resultid="7343" lane="3" heatid="8567">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="994" swimtime="00:00:28.86" resultid="7334" lane="3" heatid="8549" />
                <RESULT eventid="1414" status="DNS" swimtime="00:00:00.00" resultid="7335" lane="3" heatid="8615" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="POS" name="Poseydon" nation="RUS">
          <CONTACT email="info@dcsport.ru" name="Vera Tarasova" />
          <ATHLETES>
            <ATHLETE birthdate="1963-01-01" firstname="Vladislav" gender="M" lastname="Zagrebenko" nation="RUS" athleteid="7332">
              <RESULTS>
                <RESULT comment="World Masters Rekord" eventid="1284" points="1132" swimtime="00:00:29.47" resultid="7340" lane="4" heatid="8549" />
                <RESULT eventid="1414" status="DNS" swimtime="00:00:00.00" resultid="7341" lane="2" heatid="8615" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-SSCHVB" name="Schweiz. Schwimmvereinigung" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1991-08-15" firstname="Michael" gender="M" lastname="Greber" nation="SUI" athleteid="7449">
              <HANDICAP breast="8" free="9" medley="9" />
              <RESULTS>
                <RESULT eventid="1300" points="78" swimtime="00:00:52.04" resultid="7519" lane="1" heatid="8575" />
                <RESULT eventid="1378" points="46" swimtime="00:01:10.64" resultid="7520" lane="1" heatid="8606" />
                <RESULT eventid="1450" points="53" swimtime="00:02:11.22" resultid="7521" lane="2" heatid="8621">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="43" swimtime="00:02:34.52" resultid="7522" lane="5" heatid="8554">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-11-01" firstname="Thomas" gender="M" lastname="Wittwer" nation="SUI" athleteid="7456">
              <HANDICAP breast="4" free="6" medley="6" />
              <RESULTS>
                <RESULT eventid="1378" points="127" swimtime="00:00:57.34" resultid="7495" lane="5" heatid="8606" />
                <RESULT eventid="1284" points="98" swimtime="00:01:06.41" resultid="7493" lane="4" heatid="8545" />
                <RESULT eventid="1288" points="149" swimtime="00:02:02.59" resultid="7496" lane="2" heatid="8554">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="103" swimtime="00:02:26.40" resultid="7494" lane="3" heatid="8612">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-30" firstname="Pablo" gender="M" lastname="Gallardo" nation="SUI" athleteid="7457">
              <HANDICAP free="9" />
              <RESULTS>
                <RESULT eventid="1157" status="WDR" swimtime="00:00:00.00" resultid="7500" />
                <RESULT eventid="1300" status="WDR" swimtime="00:00:00.00" resultid="7497" />
                <RESULT eventid="1450" status="WDR" swimtime="00:00:00.00" resultid="7498" />
                <RESULT eventid="1107" status="WDR" swimtime="00:00:00.00" resultid="7499" />
                <RESULT eventid="1196" status="WDR" swimtime="00:00:00.00" resultid="7501" />
                <RESULT eventid="1292" status="WDR" swimtime="00:00:00.00" resultid="7502" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-08-31" firstname="Mirjam" gender="F" lastname="Schädler" nation="SUI" athleteid="7459">
              <HANDICAP free="6" />
              <RESULTS>
                <RESULT eventid="1286" points="19" swimtime="00:04:45.52" resultid="7510" lane="2" heatid="8550">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:14.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="22" swimtime="00:03:50.55" resultid="7509" lane="2" heatid="8616">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="18" swimtime="00:01:50.47" resultid="7508" lane="3" heatid="8569" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-05-02" firstname="Dominik" gender="M" lastname="Stäger" nation="SUI" athleteid="7472">
              <HANDICAP breast="8" free="8" medley="8" />
              <RESULTS>
                <RESULT eventid="1107" points="52" swimtime="00:04:48.07" resultid="7599" lane="5" heatid="8538">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.91" />
                    <SPLIT distance="100" swimtime="00:02:11.76" />
                    <SPLIT distance="150" swimtime="00:03:26.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="65" swimtime="00:01:03.00" resultid="7600" lane="5" heatid="8605" />
                <RESULT eventid="1288" points="56" swimtime="00:02:21.87" resultid="7601" lane="4" heatid="8553">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1450" points="48" swimtime="00:02:15.36" resultid="7598" lane="2" heatid="8620">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="61" swimtime="00:00:56.54" resultid="7597" lane="2" heatid="8574" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-13" firstname="Bruno" gender="M" lastname="Gasser" nation="SUI" athleteid="7475">
              <HANDICAP breast="10" free="10" medley="10" />
              <RESULTS>
                <RESULT eventid="1300" points="126" swimtime="00:00:46.12" resultid="7614" lane="2" heatid="8575" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-02-05" firstname="Haenni" gender="M" lastname="Walter" nation="SUI" athleteid="7476">
              <HANDICAP breast="5" free="7" medley="6" />
              <RESULTS>
                <RESULT eventid="1450" points="49" swimtime="00:02:29.56" resultid="7617" lane="5" heatid="8621">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="51" swimtime="00:01:06.00" resultid="7618" lane="6" heatid="8575" />
                <RESULT eventid="1284" points="27" swimtime="00:01:41.79" resultid="7616" lane="2" heatid="8545" />
                <RESULT eventid="1414" points="36" swimtime="00:03:26.81" resultid="7615" lane="4" heatid="8612">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="38" swimtime="00:01:25.35" resultid="7619" lane="3" heatid="8605" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-02-19" firstname="Denise" gender="F" lastname="Huser" nation="SUI" athleteid="7478">
              <HANDICAP breast="5" free="7" medley="7" />
              <RESULTS>
                <RESULT eventid="1286" points="36" swimtime="00:03:14.91" resultid="7628" lane="3" heatid="8550">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1360" points="39" swimtime="00:01:31.81" resultid="7627" lane="2" heatid="8603" />
                <RESULT eventid="1298" points="19" swimtime="00:01:39.02" resultid="7625" lane="4" heatid="8569" />
                <RESULT comment="204 - Starten vor dem Startkommando (Time: 10:40)" eventid="1432" status="DSQ" swimtime="00:03:34.16" resultid="7626" lane="3" heatid="8616">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:41.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-14" firstname="Erwin" gender="M" lastname="Dürst" nation="SUI" athleteid="8527">
              <HANDICAP breast="8" free="9" medley="9" />
              <RESULTS>
                <RESULT eventid="1300" points="211" swimtime="00:00:43.80" resultid="8528" lane="4" heatid="8575" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-WINT" name="Schwimmclub Winterthur Delfino" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1991-09-18" firstname="Stephanie" gender="F" lastname="Baumann" nation="SUI" athleteid="7450">
              <HANDICAP breast="9" free="9" medley="9" />
              <RESULTS>
                <RESULT eventid="1432" points="427" swimtime="00:01:14.12" resultid="7524" lane="3" heatid="8618">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="454" swimtime="00:00:33.30" resultid="7523" lane="3" heatid="8572" />
                <RESULT eventid="1054" points="450" swimtime="00:02:41.86" resultid="7525" lane="3" heatid="8536">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:18.21" />
                    <SPLIT distance="150" swimtime="00:02:00.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="469" swimtime="00:01:26.21" resultid="7531" lane="3" heatid="8563">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="436" swimtime="00:01:24.44" resultid="7530" lane="5" heatid="8552">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="401" swimtime="00:03:08.33" resultid="7532" lane="4" heatid="8628">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.84" />
                    <SPLIT distance="100" swimtime="00:01:30.54" />
                    <SPLIT distance="150" swimtime="00:02:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="271" swimtime="00:01:34.77" resultid="7528" lane="6" heatid="8599">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="395" swimtime="00:05:45.59" resultid="7526" lane="3" heatid="8594">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="100" swimtime="00:01:22.38" />
                    <SPLIT distance="150" swimtime="00:02:07.08" />
                    <SPLIT distance="200" swimtime="00:02:52.06" />
                    <SPLIT distance="250" swimtime="00:03:37.00" />
                    <SPLIT distance="300" swimtime="00:04:21.25" />
                    <SPLIT distance="350" swimtime="00:05:05.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1360" points="459" swimtime="00:00:38.60" resultid="7529" lane="2" heatid="8604" />
                <RESULT eventid="1396" points="344" swimtime="00:01:40.64" resultid="7527" lane="3" heatid="8610">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-04-02" firstname="Lea" gender="F" lastname="Keller" nation="SUI" athleteid="7451">
              <HANDICAP breast="5" free="6" medley="6" />
              <RESULTS>
                <RESULT eventid="1054" points="15" swimtime="00:08:14.48" resultid="7535" lane="2" heatid="8535">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:53.44" />
                    <SPLIT distance="100" swimtime="00:04:01.23" />
                    <SPLIT distance="150" swimtime="00:06:10.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="18" swimtime="00:04:01.09" resultid="7539" lane="4" heatid="8550">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:56.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="37" swimtime="00:01:37.91" resultid="7536" lane="2" heatid="8542" />
                <RESULT eventid="1298" points="11" swimtime="00:01:52.80" resultid="7533" lane="2" heatid="8569" />
                <RESULT eventid="1396" points="32" swimtime="00:03:40.45" resultid="7537" lane="4" heatid="8609">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:40.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="11" swimtime="00:04:06.26" resultid="7534" lane="4" heatid="8616">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:53.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1360" points="15" swimtime="00:01:58.79" resultid="7538" lane="5" heatid="8603" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-10-18" firstname="Giuliana" gender="F" lastname="Bavaro" nation="SUI" athleteid="7452">
              <HANDICAP breast="7" free="8" />
              <RESULTS>
                <RESULT eventid="1282" points="68" swimtime="00:01:20.09" resultid="7542" lane="3" heatid="8542" />
                <RESULT eventid="1396" points="61" swimtime="00:02:59.12" resultid="7543" lane="3" heatid="8609">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1360" points="29" swimtime="00:01:36.53" resultid="7544" lane="1" heatid="8603" />
                <RESULT eventid="1432" points="36" swimtime="00:02:48.94" resultid="7541" lane="1" heatid="8617">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.59" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="302 - Wand nicht berührt (Wende ...)" eventid="1298" status="DSQ" swimtime="00:01:20.14" resultid="7540" lane="6" heatid="8570" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-12-29" firstname="Ramona" gender="F" lastname="Loosli" nation="SUI" athleteid="7453">
              <HANDICAP breast="9" free="9" />
              <RESULTS>
                <RESULT eventid="1282" points="179" swimtime="00:00:58.17" resultid="7548" lane="5" heatid="8543" />
                <RESULT eventid="1286" points="145" swimtime="00:02:01.85" resultid="7481" lane="2" heatid="8551">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1360" points="147" swimtime="00:00:56.37" resultid="7480" lane="3" heatid="8603" />
                <RESULT eventid="1396" points="168" swimtime="00:02:07.79" resultid="7549" lane="5" heatid="8610">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="145" swimtime="00:08:02.29" resultid="7547" lane="4" heatid="8593">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.12" />
                    <SPLIT distance="100" swimtime="00:01:52.81" />
                    <SPLIT distance="150" swimtime="00:02:55.45" />
                    <SPLIT distance="200" swimtime="00:03:56.80" />
                    <SPLIT distance="250" swimtime="00:04:59.72" />
                    <SPLIT distance="300" swimtime="00:06:02.47" />
                    <SPLIT distance="350" swimtime="00:07:03.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="139" swimtime="00:00:49.41" resultid="7545" lane="6" heatid="8571" />
                <RESULT eventid="1432" points="131" swimtime="00:01:49.80" resultid="7546" lane="2" heatid="8617">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="194" swimtime="00:01:55.58" resultid="7487" lane="2" heatid="8562">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-07-14" firstname="Nicole" gender="F" lastname="Brunschwiler" nation="SUI" athleteid="7455">
              <HANDICAP breast="5" free="6" medley="6" />
              <RESULTS>
                <RESULT eventid="1282" points="15" swimtime="00:02:11.02" resultid="7490" lane="5" heatid="8542" />
                <RESULT eventid="1360" points="20" swimtime="00:01:49.59" resultid="7491" lane="2" heatid="8602" />
                <RESULT eventid="1286" points="18" swimtime="00:04:03.22" resultid="7492" lane="5" heatid="8550">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:56.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="11" swimtime="00:01:54.33" resultid="7489" lane="5" heatid="8569" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-12-04" firstname="Johannes" gender="M" lastname="Dumelin" nation="SUI" athleteid="7458">
              <HANDICAP breast="14" free="14" medley="14" />
              <RESULTS>
                <RESULT eventid="1378" points="30" swimtime="00:01:21.05" resultid="7507" lane="4" heatid="8605" />
                <RESULT eventid="1284" points="39" swimtime="00:01:22.96" resultid="7505" lane="6" heatid="8545" />
                <RESULT eventid="1450" points="29" swimtime="00:02:40.08" resultid="7504" lane="3" heatid="8620">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="40" swimtime="00:01:05.13" resultid="7503" lane="1" heatid="9290" />
                <RESULT eventid="1414" points="42" swimtime="00:02:58.60" resultid="7506" lane="2" heatid="8612">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-12-15" firstname="Sabrina" gender="F" lastname="Pfeiffer" nation="SUI" athleteid="7462">
              <HANDICAP breast="201" free="201" medley="201" />
              <RESULTS>
                <RESULT eventid="1298" points="59" swimtime="00:01:05.63" resultid="7561" lane="5" heatid="8570" />
                <RESULT eventid="1282" points="126" swimtime="00:01:05.31" resultid="7562" lane="1" heatid="8543" />
                <RESULT eventid="1360" points="78" swimtime="00:01:09.68" resultid="7564" lane="4" heatid="8602" />
                <RESULT comment="526 - Beinbewegung nicht gleichzeitig in derselben horizontalen Ebene (Time: 10:15)" eventid="1396" status="DSQ" swimtime="00:02:33.07" resultid="7563" lane="2" heatid="8609">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-12-03" firstname="Carla" gender="F" lastname="De Bortoli" nation="SUI" athleteid="7468">
              <HANDICAP breast="13" free="13" medley="13" />
              <RESULTS>
                <RESULT eventid="1396" points="360" swimtime="00:01:39.15" resultid="7586" lane="4" heatid="8610">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="348" swimtime="00:00:46.63" resultid="7585" lane="6" heatid="8544" />
                <RESULT eventid="1294" points="276" swimtime="00:01:42.85" resultid="7587" lane="4" heatid="8562">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="238" swimtime="00:06:48.79" resultid="7584" lane="2" heatid="8593">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                    <SPLIT distance="100" swimtime="00:01:35.96" />
                    <SPLIT distance="150" swimtime="00:02:28.43" />
                    <SPLIT distance="200" swimtime="00:03:22.04" />
                    <SPLIT distance="250" swimtime="00:04:16.23" />
                    <SPLIT distance="300" swimtime="00:05:10.31" />
                    <SPLIT distance="350" swimtime="00:06:02.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="219" swimtime="00:01:32.48" resultid="7583" lane="4" heatid="8617">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="270" swimtime="00:00:39.62" resultid="7582" lane="2" heatid="8571" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-11-09" firstname="Nadin" gender="F" lastname="Lüthi" nation="SUI" athleteid="7471">
              <HANDICAP breast="9" free="9" medley="9" />
              <RESULTS>
                <RESULT eventid="1302" points="125" swimtime="00:05:03.12" resultid="7594" lane="1" heatid="8582">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.19" />
                    <SPLIT distance="100" swimtime="00:02:25.04" />
                    <SPLIT distance="150" swimtime="00:03:43.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="120" swimtime="00:01:06.44" resultid="7592" lane="6" heatid="8543" />
                <RESULT eventid="1286" points="101" swimtime="00:02:17.50" resultid="7596" lane="1" heatid="8551">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" points="124" swimtime="00:02:21.33" resultid="7593" lane="1" heatid="8610">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1360" points="93" swimtime="00:01:05.58" resultid="7595" lane="4" heatid="8603" />
                <RESULT eventid="1298" points="66" swimtime="00:01:03.14" resultid="7590" lane="2" heatid="8570" />
                <RESULT eventid="1432" points="56" swimtime="00:02:25.08" resultid="7591" lane="5" heatid="8617">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-09-24" firstname="Wolf" gender="M" lastname="Schweitzer" nation="SUI" athleteid="7474">
              <HANDICAP breast="9" free="9" medley="9" />
              <RESULTS>
                <RESULT eventid="1107" points="447" swimtime="00:02:34.79" resultid="7612" lane="2" heatid="8539">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:13.55" />
                    <SPLIT distance="150" swimtime="00:01:54.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="414" swimtime="00:01:30.09" resultid="7609" lane="1" heatid="8614">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="473" swimtime="00:00:31.33" resultid="7610" lane="4" heatid="8577" />
                <RESULT eventid="1450" points="460" swimtime="00:01:09.20" resultid="7611" lane="4" heatid="8622">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="341" swimtime="00:00:38.16" resultid="7613" lane="2" heatid="8558" />
                <RESULT eventid="1284" points="336" swimtime="00:00:42.40" resultid="7608" lane="2" heatid="8546" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-05" firstname="Philipp" gender="M" lastname="Rammerstorfer" nation="SUI" athleteid="7477">
              <HANDICAP breast="2" free="3" />
              <RESULTS>
                <RESULT eventid="1288" points="15" swimtime="00:03:36.23" resultid="7624" lane="6" heatid="8554">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:45.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1378" points="14" swimtime="00:01:44.37" resultid="7623" lane="2" heatid="8605" />
                <RESULT eventid="1284" points="4" swimtime="00:02:46.42" resultid="7622" lane="1" heatid="8545" />
                <RESULT eventid="1450" points="10" swimtime="00:03:45.58" resultid="7621" lane="4" heatid="8620">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:48.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="12" swimtime="00:01:35.44" resultid="7620" lane="3" heatid="8574" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-CHUR" name="Schwimmclub Chur" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1994-04-26" firstname="Madlaina" gender="F" lastname="Gaudenz" nation="SUI" athleteid="7454">
              <HANDICAP breast="8" free="10" medley="9" />
              <RESULTS>
                <RESULT eventid="1290" points="310" swimtime="00:00:40.74" resultid="8723" lane="5" heatid="8557" />
                <RESULT eventid="1294" points="318" swimtime="00:01:38.08" resultid="7488" lane="3" heatid="8562">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="350" swimtime="00:01:30.90" resultid="7486" lane="6" heatid="8552">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="315" swimtime="00:00:37.61" resultid="7482" lane="1" heatid="8572" />
                <RESULT eventid="1432" points="341" swimtime="00:01:19.86" resultid="7483" lane="1" heatid="8618">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1054" points="391" swimtime="00:02:49.57" resultid="7484" lane="1" heatid="8536">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:21.18" />
                    <SPLIT distance="150" swimtime="00:02:06.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="353" swimtime="00:05:58.74" resultid="7485" lane="5" heatid="8594">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                    <SPLIT distance="100" swimtime="00:01:25.30" />
                    <SPLIT distance="150" swimtime="00:02:10.97" />
                    <SPLIT distance="200" swimtime="00:02:56.42" />
                    <SPLIT distance="250" swimtime="00:03:42.13" />
                    <SPLIT distance="300" swimtime="00:04:27.68" />
                    <SPLIT distance="350" swimtime="00:05:13.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1360" points="338" swimtime="00:00:42.73" resultid="9856" lane="3" heatid="8602" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-GER" name="Behindertenschwimmer Germany" nation="GER">
          <ATHLETES>
            <ATHLETE birthdate="1962-03-08" firstname="Markus" gender="M" lastname="Schnitzer" nation="GER" athleteid="7460">
              <HANDICAP free="10" medley="10" />
              <RESULTS>
                <RESULT eventid="1378" points="390" swimtime="00:00:39.50" resultid="7514" lane="6" heatid="8607" />
                <RESULT eventid="1107" points="407" swimtime="00:02:45.37" resultid="7511" lane="4" heatid="8539">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:19.89" />
                    <SPLIT distance="150" swimtime="00:02:03.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="321" swimtime="00:13:22.98" resultid="7513" lane="5" heatid="8589">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                    <SPLIT distance="100" swimtime="00:01:31.77" />
                    <SPLIT distance="150" swimtime="00:02:19.63" />
                    <SPLIT distance="200" swimtime="00:03:08.01" />
                    <SPLIT distance="250" swimtime="00:03:57.13" />
                    <SPLIT distance="300" swimtime="00:04:46.96" />
                    <SPLIT distance="350" swimtime="00:05:37.70" />
                    <SPLIT distance="400" swimtime="00:06:29.24" />
                    <SPLIT distance="450" swimtime="00:07:20.71" />
                    <SPLIT distance="500" swimtime="00:08:12.70" />
                    <SPLIT distance="550" swimtime="00:09:04.81" />
                    <SPLIT distance="600" swimtime="00:09:56.95" />
                    <SPLIT distance="650" swimtime="00:10:49.07" />
                    <SPLIT distance="700" swimtime="00:11:40.84" />
                    <SPLIT distance="750" swimtime="00:12:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="394" swimtime="00:05:58.20" resultid="7512" lane="4" heatid="8596">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                    <SPLIT distance="100" swimtime="00:01:24.71" />
                    <SPLIT distance="150" swimtime="00:02:09.42" />
                    <SPLIT distance="200" swimtime="00:02:55.53" />
                    <SPLIT distance="250" swimtime="00:03:40.86" />
                    <SPLIT distance="300" swimtime="00:04:26.74" />
                    <SPLIT distance="350" swimtime="00:05:12.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="440" swimtime="00:01:25.55" resultid="7550" lane="1" heatid="8555">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="286" swimtime="00:01:36.47" resultid="7551" lane="5" heatid="8565">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1486" points="490" swimtime="00:02:58.70" resultid="9092" lane="2" heatid="8626">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                    <SPLIT distance="100" swimtime="00:01:27.31" />
                    <SPLIT distance="150" swimtime="00:02:13.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1522" points="317" swimtime="00:03:25.07" resultid="9095" lane="6" heatid="8630">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.47" />
                    <SPLIT distance="100" swimtime="00:01:43.52" />
                    <SPLIT distance="150" swimtime="00:02:41.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-SKWORB" name="Schwimmklub Worb" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1978-02-12" firstname="Chantal" gender="F" lastname="Cavin" nation="SUI" athleteid="7461">
              <HANDICAP breast="11" free="11" medley="11" />
              <RESULTS>
                <RESULT eventid="1290" points="402" swimtime="00:00:39.05" resultid="7558" lane="2" heatid="8557" />
                <RESULT eventid="1324" points="259" swimtime="00:01:40.24" resultid="7559" lane="1" heatid="8599">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="350" swimtime="00:01:32.21" resultid="7560" lane="2" heatid="8563">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="315" swimtime="00:00:48.88" resultid="7556" lane="1" heatid="8544" />
                <RESULT eventid="1298" points="529" swimtime="00:00:32.85" resultid="7552" lane="5" heatid="8573" />
                <RESULT eventid="1432" points="456" swimtime="00:01:15.43" resultid="7553" lane="6" heatid="8619">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Behinderten Weltrekord S11 (blind)" eventid="1054" points="493" swimtime="00:02:38.59" resultid="7554" lane="6" heatid="8537">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:16.59" />
                    <SPLIT distance="150" swimtime="00:01:59.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="462" swimtime="00:05:46.72" resultid="7555" lane="2" heatid="8594">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                    <SPLIT distance="100" swimtime="00:01:24.89" />
                    <SPLIT distance="150" swimtime="00:02:08.88" />
                    <SPLIT distance="200" swimtime="00:02:52.91" />
                    <SPLIT distance="250" swimtime="00:03:37.16" />
                    <SPLIT distance="300" swimtime="00:04:21.88" />
                    <SPLIT distance="350" swimtime="00:05:06.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1396" status="WDR" swimtime="00:00:00.00" resultid="7557" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-SVK" name="Schwimmverein Kriens" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1990-05-08" firstname="Andrea" gender="F" lastname="Seiler" nation="SUI" athleteid="7463">
              <HANDICAP breast="9" free="9" medley="9" />
              <RESULTS>
                <RESULT eventid="1432" points="372" swimtime="00:01:17.60" resultid="7566" lane="6" heatid="8618">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1360" points="383" swimtime="00:00:41.01" resultid="7568" lane="1" heatid="8604" />
                <RESULT eventid="1286" points="338" swimtime="00:01:31.95" resultid="7569" lane="1" heatid="8552">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1468" points="320" swimtime="00:03:18.24" resultid="7570" lane="2" heatid="8625">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:35.85" />
                    <SPLIT distance="150" swimtime="00:02:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="407" swimtime="00:01:30.34" resultid="7571" lane="1" heatid="8563">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="372" swimtime="00:00:35.60" resultid="7565" lane="5" heatid="8572" />
                <RESULT eventid="1054" points="365" swimtime="00:02:53.47" resultid="7567" lane="6" heatid="8536">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                    <SPLIT distance="150" swimtime="00:02:07.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-BSGZ" name="Behindertensportgruppe Zimmerberg" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1984-11-23" firstname="Philipp" gender="M" lastname="Leuzinger" nation="SUI" athleteid="7464">
              <HANDICAP breast="9" free="9" medley="9" />
              <RESULTS>
                <RESULT eventid="1107" points="61" swimtime="00:04:39.86" resultid="7573" lane="4" heatid="8538">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.73" />
                    <SPLIT distance="100" swimtime="00:02:10.43" />
                    <SPLIT distance="150" swimtime="00:03:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="203 - Bewegen vor dem Startkommando" eventid="1300" status="DSQ" swimtime="00:00:51.41" resultid="7572" lane="5" heatid="8575" />
                <RESULT comment="Schwimmen auf Bauchlage - Aufgegeben" eventid="1288" status="DSQ" swimtime="00:00:00.00" resultid="7574" lane="2" heatid="8553">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-08-07" firstname="Matthias" gender="M" lastname="Rusterholz" nation="SUI" athleteid="7465">
              <HANDICAP breast="9" free="9" medley="9" />
              <RESULTS>
                <RESULT eventid="1288" points="77" swimtime="00:02:11.88" resultid="7576" lane="3" heatid="8553">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="128" swimtime="00:00:45.07" resultid="7575" lane="6" heatid="8574" />
                <RESULT eventid="1296" status="WDR" swimtime="00:00:00.00" resultid="7577" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-02-08" firstname="Nicole" gender="F" lastname="Odermatt" nation="SUI" athleteid="7466">
              <HANDICAP breast="7" free="7" medley="7" />
              <RESULTS>
                <RESULT eventid="1286" points="97" swimtime="00:02:19.20" resultid="7579" lane="5" heatid="8551">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="91" swimtime="00:00:56.78" resultid="7578" lane="3" heatid="8570" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-12-02" firstname="Cécile" gender="F" lastname="Bucher" nation="SUI" athleteid="7467">
              <HANDICAP breast="7" free="8" medley="8" />
              <RESULTS>
                <RESULT eventid="1286" points="75" swimtime="00:02:31.47" resultid="7581" lane="6" heatid="8551">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="23" swimtime="00:01:28.96" resultid="7580" lane="1" heatid="8570" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Basil" gender="M" lastname="Dias" nation="SUI" athleteid="7469">
              <HANDICAP breast="6" free="7" medley="7" />
              <RESULTS>
                <RESULT eventid="1300" points="3" swimtime="00:02:21.39" resultid="7588" lane="4" heatid="8574" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-10-25" firstname="Svonislav" gender="M" lastname="Jankovic" nation="SUI" athleteid="7470">
              <HANDICAP breast="201" free="201" medley="201" />
              <RESULTS>
                <RESULT eventid="1300" points="25" swimtime="00:01:15.88" resultid="7589" lane="5" heatid="8574" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-LIMM" name="SV Limmat Sharks" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1974-07-03" firstname="Reto" gender="M" lastname="Thurnherr" nation="SUI" athleteid="7473">
              <HANDICAP breast="8" free="8" medley="8" />
              <RESULTS>
                <RESULT eventid="1157" points="272" swimtime="00:06:18.54" resultid="7605" lane="5" heatid="8597">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.63" />
                    <SPLIT distance="100" swimtime="00:01:26.56" />
                    <SPLIT distance="150" swimtime="00:02:14.00" />
                    <SPLIT distance="200" swimtime="00:03:02.41" />
                    <SPLIT distance="250" swimtime="00:03:51.80" />
                    <SPLIT distance="300" swimtime="00:04:40.96" />
                    <SPLIT distance="350" swimtime="00:05:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1450" points="241" swimtime="00:01:22.61" resultid="7603" lane="6" heatid="8622">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="228" swimtime="00:00:41.15" resultid="7606" lane="3" heatid="8558" />
                <RESULT eventid="1107" points="271" swimtime="00:02:59.44" resultid="7604" lane="6" heatid="8539">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                    <SPLIT distance="100" swimtime="00:01:23.81" />
                    <SPLIT distance="150" swimtime="00:02:11.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="233" swimtime="00:00:37.61" resultid="7602" lane="1" heatid="8576" />
                <RESULT eventid="1296" points="182" swimtime="00:01:43.03" resultid="7607" lane="6" heatid="8565">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-BSGO" name="BSG Obwalden" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1985-08-17" firstname="Corinne" gender="F" lastname="Gasser" nation="SUI" athleteid="7479">
              <HANDICAP breast="14" free="14" medley="14" />
              <RESULTS>
                <RESULT eventid="1298" points="94" swimtime="00:00:56.22" resultid="7629" lane="4" heatid="8570" />
                <RESULT comment="303 - Nicht mit beiden Händen gleich-zeitig angeschlagen (Wende  ...)" eventid="1282" status="DSQ" swimtime="00:01:05.16" resultid="7630" lane="4" heatid="8542" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SSG" name="SSG Saar MR" nation="GER">
          <CONTACT city="Friedrichsthal" country="DE" email="AnneSchmitt-SSG@web.de" name="Anne Schmitt" phone="0171 15 74 103" street="Ludwigstrasse 10" zip="66299" />
          <ATHLETES>
            <ATHLETE birthdate="1940-01-01" firstname="Hermann" gender="M" lastname="Sittner" nation="GER" license="93461" athleteid="7665">
              <RESULTS>
                <RESULT eventid="1304" points="370" swimtime="00:04:16.93" resultid="7667" lane="5" heatid="8583">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.30" />
                    <SPLIT distance="100" swimtime="00:02:01.83" />
                    <SPLIT distance="150" swimtime="00:03:10.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="360" swimtime="00:00:50.86" resultid="7666" lane="3" heatid="8545" />
                <RESULT eventid="1414" points="376" swimtime="00:01:52.82" resultid="7668" lane="5" heatid="8613">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TV 1872" name="TV 1872 Saarlouis" nation="FRA">
          <CONTACT city="Creutzwald" country="FR" name="Kurt Mayer" street="60 rue du Maréchal Ney" zip="57150" />
          <ATHLETES>
            <ATHLETE birthdate="1927-01-01" firstname="Kurt" gender="M" lastname="Mayer" nation="FRA" license="135080" athleteid="7670">
              <RESULTS>
                <RESULT eventid="1378" points="136" swimtime="00:01:19.55" resultid="7673" lane="6" heatid="8606" />
                <RESULT eventid="1486" points="158" swimtime="00:06:19.44" resultid="7674" lane="4" heatid="8626">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.39" />
                    <SPLIT distance="100" swimtime="00:03:08.10" />
                    <SPLIT distance="150" swimtime="00:04:48.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="144" swimtime="00:01:25.79" resultid="7671" lane="5" heatid="8545" />
                <RESULT eventid="1288" points="158" swimtime="00:02:51.99" resultid="7672" lane="1" heatid="8554">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GEN" name="Genève Natation 1885" nation="SUI" region="RSR">
          <CONTACT city="Genève 26" email="info@geneve-natation-1885.ch" fax="022/301.36.96" name="Secrétariat" phone="022/342.19.72" street="Piscine des Vernets" street2="Velardo Patricia" zip="CH-1211" />
          <ATHLETES>
            <ATHLETE birthdate="1959-07-18" firstname="Robert" gender="M" lastname="Alderton" nation="GBR" athleteid="7812">
              <RESULTS>
                <RESULT eventid="1378" status="DNS" swimtime="00:00:00.00" resultid="7816" lane="4" heatid="8608" />
                <RESULT eventid="1296" status="DNS" swimtime="00:00:00.00" resultid="7815" lane="3" heatid="8566" />
                <RESULT eventid="1486" status="DNS" swimtime="00:00:00.00" resultid="7817" lane="4" heatid="8627" />
                <RESULT eventid="1284" status="DNS" swimtime="00:00:00.00" resultid="7813" lane="5" heatid="8548" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="7814" lane="3" heatid="8556" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-12-12" firstname="Jonathan" gender="M" lastname="Banville" nation="CAN" license="15297" athleteid="7818">
              <RESULTS>
                <RESULT eventid="1414" points="852" swimtime="00:01:06.76" resultid="7822" lane="4" heatid="8615">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1522" points="772" swimtime="00:02:16.71" resultid="7823" lane="3" heatid="8631">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="100" swimtime="00:01:06.31" />
                    <SPLIT distance="150" swimtime="00:01:45.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="828" swimtime="00:02:30.96" resultid="7821" lane="3" heatid="8584">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:12.69" />
                    <SPLIT distance="150" swimtime="00:01:51.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="769" swimtime="00:01:03.74" resultid="7820" lane="4" heatid="8567">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="750" swimtime="00:00:31.70" resultid="7819" lane="2" heatid="8549" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-08-06" firstname="Andreas" gender="M" lastname="Herty" nation="GER" license="18212" athleteid="7836">
              <RESULTS>
                <RESULT eventid="1378" points="413" swimtime="00:00:35.06" resultid="7839" lane="5" heatid="8608" />
                <RESULT eventid="1486" points="407" swimtime="00:02:50.52" resultid="7840" lane="6" heatid="8627">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:22.16" />
                    <SPLIT distance="150" swimtime="00:02:07.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="418" swimtime="00:01:17.91" resultid="7838" lane="4" heatid="8566">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="388" swimtime="00:01:17.64" resultid="7837" lane="5" heatid="8556">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-19" firstname="Daniela" gender="F" lastname="Menegon" nation="ITA" license="22084" athleteid="7847">
              <RESULTS>
                <RESULT eventid="1054" points="665" swimtime="00:02:23.54" resultid="7848" lane="2" heatid="8537">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:10.32" />
                    <SPLIT distance="150" swimtime="00:01:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="587" swimtime="00:00:31.74" resultid="7849" lane="2" heatid="8573" />
                <RESULT eventid="1177" points="721" swimtime="00:10:30.27" resultid="7850" lane="2" heatid="8588">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="150" swimtime="00:01:51.22" />
                    <SPLIT distance="200" swimtime="00:02:30.04" />
                    <SPLIT distance="250" swimtime="00:03:08.74" />
                    <SPLIT distance="300" swimtime="00:03:47.73" />
                    <SPLIT distance="350" swimtime="00:04:27.48" />
                    <SPLIT distance="400" swimtime="00:05:07.22" />
                    <SPLIT distance="450" swimtime="00:05:47.43" />
                    <SPLIT distance="500" swimtime="00:06:27.77" />
                    <SPLIT distance="550" swimtime="00:07:08.16" />
                    <SPLIT distance="600" swimtime="00:07:48.53" />
                    <SPLIT distance="650" swimtime="00:08:29.17" />
                    <SPLIT distance="700" swimtime="00:09:09.86" />
                    <SPLIT distance="750" swimtime="00:09:50.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="658" swimtime="00:05:08.22" resultid="7851" lane="5" heatid="8595">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                    <SPLIT distance="150" swimtime="00:01:51.34" />
                    <SPLIT distance="200" swimtime="00:02:30.46" />
                    <SPLIT distance="250" swimtime="00:03:10.01" />
                    <SPLIT distance="300" swimtime="00:03:49.45" />
                    <SPLIT distance="350" swimtime="00:04:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="623" swimtime="00:01:07.96" resultid="7852" lane="2" heatid="8619">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1504" points="536" swimtime="00:02:55.90" resultid="7853" lane="3" heatid="8628">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:01:26.52" />
                    <SPLIT distance="150" swimtime="00:02:15.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-02-21" firstname="Simon" gender="M" lastname="Pagin" nation="SUI" license="16719" athleteid="7854">
              <RESULTS>
                <RESULT eventid="1284" points="444" swimtime="00:00:42.19" resultid="7857" lane="4" heatid="8546" />
                <RESULT eventid="1342" points="390" swimtime="00:01:26.41" resultid="7856" lane="3" heatid="8600">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="525" swimtime="00:00:34.37" resultid="7858" lane="1" heatid="8560" />
                <RESULT eventid="1300" points="563" swimtime="00:00:30.72" resultid="7855" lane="3" heatid="8577" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="VN" name="Vevey Natation" nation="SUI">
          <CONTACT email="cmswisschris@gmail.com" name="Morgan Chris" />
          <ATHLETES>
            <ATHLETE birthdate="1969-01-01" firstname="Chris" gender="M" lastname="Morgan" nation="SUI" athleteid="7868">
              <RESULTS>
                <RESULT eventid="1292" points="938" swimtime="00:00:27.23" resultid="7870" lane="4" heatid="8561" />
                <RESULT eventid="1300" points="837" swimtime="00:00:25.91" resultid="7871" lane="5" heatid="8581" />
                <RESULT eventid="1196" points="556" swimtime="00:10:29.35" resultid="8750" lane="6" heatid="8589">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="100" swimtime="00:01:08.74" />
                    <SPLIT distance="150" swimtime="00:01:46.93" />
                    <SPLIT distance="200" swimtime="00:02:25.60" />
                    <SPLIT distance="250" swimtime="00:03:04.19" />
                    <SPLIT distance="300" swimtime="00:03:43.91" />
                    <SPLIT distance="350" swimtime="00:04:24.26" />
                    <SPLIT distance="400" swimtime="00:05:04.71" />
                    <SPLIT distance="450" swimtime="00:05:44.96" />
                    <SPLIT distance="500" swimtime="00:06:26.42" />
                    <SPLIT distance="550" swimtime="00:07:07.53" />
                    <SPLIT distance="600" swimtime="00:07:48.68" />
                    <SPLIT distance="650" swimtime="00:08:29.32" />
                    <SPLIT distance="700" swimtime="00:09:10.13" />
                    <SPLIT distance="750" swimtime="00:09:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="737" swimtime="00:02:11.03" resultid="7869" lane="5" heatid="8540">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="100" swimtime="00:01:02.91" />
                    <SPLIT distance="150" swimtime="00:01:37.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ASA" name="ASA Nuoto Cinisello ASD" nation="ITA">
          <CONTACT city="Cinisello Balsamo MI" country="IT" email="max.cassaghi@alice.it" name="Massimo Cassaghi" phone="0039 349 2259313" street="Via Vittorio Veneto 17" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Massimo" gender="M" lastname="Cassaghi" nation="ITA" license="LOM 035429" athleteid="7875">
              <RESULTS>
                <RESULT eventid="1378" points="714" swimtime="00:00:31.34" resultid="7876" lane="2" heatid="8608" />
                <RESULT eventid="1450" points="778" swimtime="00:00:58.06" resultid="7877" lane="5" heatid="8624">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOSIR" name="Mosir" nation="POL" shortname="MOSIR">
          <ATHLETES>
            <ATHLETE birthdate="1945-01-01" firstname="Jozef" gender="M" lastname="Rozalski" nation="POL" athleteid="7209">
              <RESULTS>
                <RESULT eventid="1304" points="604" swimtime="00:03:28.75" resultid="7224" lane="4" heatid="8583">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="100" swimtime="00:01:41.44" />
                    <SPLIT distance="150" swimtime="00:02:38.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="607" swimtime="00:01:22.73" resultid="7226" lane="2" heatid="8600">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="618" swimtime="00:01:32.70" resultid="7227" lane="6" heatid="8614">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="747" swimtime="00:00:30.07" resultid="7223" lane="1" heatid="8577" />
                <RESULT eventid="1522" points="622" swimtime="00:03:08.74" resultid="7229" lane="1" heatid="8630">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:01:32.62" />
                    <SPLIT distance="150" swimtime="00:02:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1450" points="681" swimtime="00:01:10.87" resultid="7228" lane="1" heatid="8622">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="582" swimtime="00:01:26.09" resultid="7222" lane="6" heatid="8566">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="577" swimtime="00:00:41.15" resultid="7220" lane="1" heatid="8546" />
                <RESULT eventid="1292" points="751" swimtime="00:00:33.41" resultid="7221" lane="3" heatid="8559" />
                <RESULT eventid="1107" points="641" swimtime="00:02:43.76" resultid="7219" lane="1" heatid="8539">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                    <SPLIT distance="100" swimtime="00:01:18.94" />
                    <SPLIT distance="150" swimtime="00:02:03.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="576" swimtime="00:05:54.65" resultid="7225" lane="2" heatid="8596">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:23.62" />
                    <SPLIT distance="150" swimtime="00:02:09.58" />
                    <SPLIT distance="200" swimtime="00:02:55.20" />
                    <SPLIT distance="250" swimtime="00:03:40.86" />
                    <SPLIT distance="300" swimtime="00:04:26.05" />
                    <SPLIT distance="350" swimtime="00:05:10.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="UNATTACHED" name="unattached">
          <OFFICIALS>
            <OFFICIAL officialid="7660" firstname="Christian" gender="M" grade="Schiiedsrichter A" lastname="Fahrni" />
          </OFFICIALS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
