<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 2007" registration="Splash Software" version="DEBUG Build">
    <CONTACT name="GeoLogix AG" street="Muristrasse 60" city="Bern" zip="3006" country="CH" phone="+41 31 356 80 56" fax="+41 31 356 80 81" email="info@splash-software.ch" internet="http://www.splash-software.ch" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Nottwil" name="Schweizerische Masters Meisterschaften" name.en="Swiss Masters Championships" course="SCM" deadline="2009-09-07" nation="SUI" organizer="Schwimmverein Emmen" state="LU" timing="AUTOMATIC" type="SUI.MCS">
      <AGEDATE value="2009-09-27" type="YEAR" />
      <POOL name="Hallenbad -- Schweiz. Paraplegikerzentrum" lanemin="1" lanemax="6" />
      <POINTTABLE pointtableid="1008" name="DSV Master Performance Table" version="2004" />
      <CONTACT city="Hildisrieden" email="info@sv-emmen.ch" internet="www.sv-emmen.ch" name="Daniel Kuratli" street="Länzeweid 33b" zip="6024" />
      <SESSIONS>
        <SESSION date="2009-09-26" daytime="13:00" name="Samstag -- Einzelwettkämpfe" number="1" officialmeeting="12:15" teamleadermeeting="12:00" warmupfrom="11:30" warmupuntil="12:45">
          <EVENTS>
            <EVENT eventid="1054" daytime="13:00" gender="F" number="1" order="1" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1070" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="1056" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="1057" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="1058" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1059" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1060" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="1061" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="1062" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="1063" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1064" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1065" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1066" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1067" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1068" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1069" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="6581" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="6582" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="6580" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="6583" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="10537" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8535" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8536" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8537" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="13:15" gender="M" number="2" order="2" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11154" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11155" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11156" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11157" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11158" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11159" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11160" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11161" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11162" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11163" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11164" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11165" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11166" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11167" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11168" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11169" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11170" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11171" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11172" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11173" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8538" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8539" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8540" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8541" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1282" daytime="13:35" gender="F" number="3" order="3" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11174" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11175" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11176" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11177" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11178" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11179" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11180" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11181" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11182" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11183" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11184" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11185" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11186" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11187" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11188" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11189" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11190" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11191" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11192" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11193" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8542" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8543" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8544" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1284" daytime="13:45" gender="M" number="4" order="4" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11194" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11195" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11196" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11197" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11198" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11199" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11200" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11201" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11202" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11203" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11204" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11205" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11206" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11207" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11208" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11209" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11210" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11211" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11212" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11213" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8545" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8546" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8547" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8548" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8549" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1286" daytime="13:55" gender="F" number="5" order="5" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11214" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11215" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11216" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11217" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11218" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11219" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11220" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11221" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11222" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11223" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11224" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11225" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11226" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11227" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11228" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11229" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11230" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11231" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11232" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11233" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8550" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8551" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8552" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1288" daytime="14:10" gender="M" number="6" order="6" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11234" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11235" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11236" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11237" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11238" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11239" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11240" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11241" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11242" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11243" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11244" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11245" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11246" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11247" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11248" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11249" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11250" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11251" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11252" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11253" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8553" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8554" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8555" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8556" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1290" daytime="14:25" gender="F" number="7" order="7" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11254" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11255" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11256" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11257" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11258" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11259" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11260" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11261" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11262" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11263" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11264" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11265" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11266" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11267" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11268" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11269" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11270" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11271" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11272" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11273" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8557" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1292" daytime="14:25" gender="M" number="8" order="8" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11274" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11275" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11276" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11277" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11278" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11279" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11280" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11281" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11282" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11283" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11284" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11285" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11286" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11287" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11288" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11289" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11290" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11291" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11292" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11293" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8558" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8559" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8560" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8561" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1294" daytime="14:35" gender="F" number="9" order="9" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11294" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11295" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11296" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11297" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11298" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11299" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11300" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11301" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11302" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11303" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11304" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11305" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11306" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11307" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11308" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11309" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11310" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11311" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11312" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11313" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8562" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8563" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8564" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1296" daytime="14:45" gender="M" number="10" order="10" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11314" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11315" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11316" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11317" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11318" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11319" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11320" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11321" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11322" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11323" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11324" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11325" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11326" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11327" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11328" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11329" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11330" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11331" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11332" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11333" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8565" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8566" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8567" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1298" daytime="14:55" gender="F" number="11" order="11" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11334" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11335" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11336" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11337" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11338" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11339" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11340" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11341" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11342" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11343" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11344" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11345" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11346" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11347" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11348" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11349" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11350" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11351" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11352" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11353" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8569" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8570" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8571" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8572" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8573" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1300" daytime="15:10" gender="M" number="12" order="12" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11354" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11355" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11356" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11357" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11358" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11359" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11360" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11361" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11362" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11363" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11364" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11365" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11366" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11367" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11368" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11369" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11370" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11371" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11372" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11373" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8574" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8575" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8576" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8577" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8578" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8579" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8580" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8581" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="9290" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1302" daytime="15:25" gender="F" number="13" order="13" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11374" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11375" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11376" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11377" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11378" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11379" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11380" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11381" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11382" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11383" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11384" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11385" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11386" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11387" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11388" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11389" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11390" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11391" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11392" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11393" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8582" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1304" daytime="15:35" gender="M" number="14" order="14" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11394" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11395" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11396" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11397" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11398" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11399" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11400" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11401" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11402" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11403" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11404" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11405" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11406" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11407" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11408" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11409" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11410" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11411" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11412" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11413" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8583" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8584" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-26" daytime="15:50" name="Samstag -- Staffeln" number="2">
          <EVENTS>
            <EVENT eventid="1175" daytime="15:50" gender="X" number="15" order="8" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="2000" />
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <HEATS>
                <HEAT heatid="8585" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-26" daytime="16:00" name="Samstag -- 800 m" number="3">
          <EVENTS>
            <EVENT eventid="1177" daytime="16:00" gender="F" number="16" order="8" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11414" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11415" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11416" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11417" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11418" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11419" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11420" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11421" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11422" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11423" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11424" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11425" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11426" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11427" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11428" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11429" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11430" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11431" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11432" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11433" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8587" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8588" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1196" daytime="16:35" gender="M" number="17" order="9" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11434" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11435" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11436" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11437" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11438" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11439" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11440" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11441" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11442" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11443" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11444" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11445" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11446" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11447" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11448" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11449" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11450" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11451" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11452" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11453" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8589" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8590" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="9736" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-27" name="Samstag  -- 1500m" number="4">
          <EVENTS>
            <EVENT eventid="7347" number="18" order="2" preveventid="-1" round="TIM">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="8592" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-27" daytime="09:00" name="Sonntag -- Einzelwettkämpfe" number="7" officialmeeting="08:30" teamleadermeeting="08:15" warmupfrom="08:00" warmupuntil="08:45">
          <EVENTS>
            <EVENT eventid="1072" daytime="09:00" gender="F" number="19" order="2" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11454" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11455" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11456" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11457" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11458" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11459" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11460" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11461" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11462" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11463" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11464" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11465" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11466" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11467" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11468" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11469" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11470" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11471" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11472" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11473" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8593" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8594" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8595" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1157" daytime="09:25" gender="M" number="20" order="3" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11474" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11475" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11476" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11477" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11478" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11479" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11480" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11481" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11482" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11483" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11484" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11485" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11486" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11487" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11488" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11489" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11490" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11491" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11492" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11493" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8596" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8597" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8598" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" daytime="09:55" gender="F" number="21" order="4" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10902" agemax="17" agemin="-1" />
                <AGEGROUP agegroupid="10903" agemax="24" agemin="18" />
                <AGEGROUP agegroupid="10904" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="10905" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="10906" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="10907" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="10908" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="10909" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="10910" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="10911" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="10912" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10913" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10914" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10915" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="10916" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="10917" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="10918" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="10919" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="10920" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="10921" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="10922" agemax="-1" agemin="-1" name="Klassierung nach Zeit" type="MASTERS" />
                <AGEGROUP agegroupid="11494" agemax="-1" agemin="-1" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8599" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1342" daytime="10:00" gender="M" number="22" order="5" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11495" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11496" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11497" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11498" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11499" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11500" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11501" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11502" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11503" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11504" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11505" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11506" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11507" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11508" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11509" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11510" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11511" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11512" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11513" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11514" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8600" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8601" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1360" daytime="10:10" gender="F" number="23" order="6" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11515" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11516" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11517" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11518" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11519" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11520" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11521" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11522" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11523" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11524" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11525" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11526" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11527" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11528" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11529" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11530" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11531" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11532" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11533" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11534" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8602" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8603" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8604" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1378" daytime="10:20" gender="M" number="24" order="7" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11535" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11536" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11537" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11538" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11539" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11540" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11541" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11542" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11543" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11544" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11545" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11546" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11547" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11548" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11549" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11550" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11551" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11552" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11553" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11554" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8605" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8606" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8607" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8608" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1396" daytime="10:30" gender="F" number="25" order="8" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11555" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11556" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11557" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11558" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11559" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11560" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11561" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11562" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11563" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11564" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11565" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11566" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11567" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11568" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11569" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11570" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11571" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11572" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11573" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11574" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8609" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8610" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8611" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1414" daytime="10:40" gender="M" number="26" order="9" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11575" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11576" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11577" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11578" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11579" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11580" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11581" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11582" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11583" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11584" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11585" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11586" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11587" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11588" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11589" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11590" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11591" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11592" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11593" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11594" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8612" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8613" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8614" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8615" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1432" daytime="10:55" gender="F" number="27" order="10" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11595" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11596" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11597" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11598" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11599" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11600" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11601" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11602" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11603" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11604" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11605" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11606" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11607" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11608" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11609" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11610" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11611" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11612" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11613" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11614" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8616" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8617" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8618" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8619" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1450" daytime="11:10" gender="M" number="28" order="11" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11615" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11616" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11617" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11618" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11619" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11620" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11621" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11622" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11623" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11624" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11625" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11626" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11627" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11628" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11629" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11630" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11631" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11632" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11633" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11634" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8620" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8621" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8622" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8623" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8624" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1468" daytime="11:25" gender="F" number="29" order="12" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11635" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11636" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11637" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11638" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11639" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11640" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11641" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11642" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11643" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11644" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11645" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11646" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11647" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11648" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11649" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11650" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11651" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11652" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11653" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11654" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8625" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1486" daytime="11:30" gender="M" number="30" order="13" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11655" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11656" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11657" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11658" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11659" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11660" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11661" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11662" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11663" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11664" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11665" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11666" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11667" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11668" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11669" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11670" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11671" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11672" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11673" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11674" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8626" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8627" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1504" daytime="11:45" gender="F" number="31" order="14" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11675" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11676" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11677" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11678" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11679" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11680" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11681" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11682" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11683" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11684" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11685" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11686" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11687" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11688" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11689" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11690" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11691" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11692" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11693" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11694" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8628" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8629" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1522" daytime="11:55" gender="M" number="32" order="15" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="1200" />
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11695" agemax="24" agemin="19" name="Pre-Masters" />
                <AGEGROUP agegroupid="11696" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="11697" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="11698" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="11699" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="11700" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="11701" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="11702" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="11703" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="11704" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="11705" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="11706" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="11707" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="11708" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="11709" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="11710" agemax="18" agemin="-1" name="SSCHVB -- Jugend S1 - S15" />
                <AGEGROUP agegroupid="11711" agemax="18" agemin="-1" name="SSCHVB -- Jugend AB" />
                <AGEGROUP agegroupid="11712" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene S1 - S15" />
                <AGEGROUP agegroupid="11713" agemax="-1" agemin="19" name="SSCHVB -- Erwachsene AB" />
                <AGEGROUP agegroupid="11714" agemax="-1" agemin="-1" name="Klassierung nach Zeit" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8630" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8631" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-27" daytime="12:10" name="Sonntag -- Staffeln" number="8">
          <EVENTS>
            <EVENT eventid="1540" daytime="12:10" gender="X" number="33" order="17" preveventid="-1" round="TIM">
              <FEE currency="CHF" value="2000" />
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT heatid="8633" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="7660" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2009-09-27" name="Staffeln der Behinderten" number="9">
          <EVENTS>
            <EVENT eventid="7349" number="35" order="21" preveventid="-1" round="TIM">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7357" agemax="-1" agemin="-1" name="Behinderte (Klasse 20)" />
                <AGEGROUP agegroupid="7350" agemax="-1" agemin="-1" name="Behinderte (Klasse 34)" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="11716" number="34" order="20" preveventid="-1" round="TIM">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11718" agemax="-1" agemin="-1" name="Behinderte (Klasse 20)" />
                <AGEGROUP agegroupid="11719" agemax="-1" agemin="-1" name="Behinderte (Klasse 34)" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="WAED" name="Schwimmverein Wädenswil" nation="SUI" region="RZO">
          <CONTACT city="Wädenswil" name="Truttmann Otto" phone="044 780 75 06" street="Freiherrenstrasse 4" zip="8820" />
          <ATHLETES>
            <ATHLETE birthdate="1954-01-12" firstname="Ales" gender="M" lastname="Vrana" nation="SUI" license="19251" athleteid="6774">
              <ENTRIES>
                <ENTRY entrytime="00:01:22.55" eventid="1414" lane="5" heatid="8614">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.83" eventid="1284" lane="4" heatid="8547">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:03:02.97" eventid="1304" lane="1" heatid="8584">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SV 01" name="Mainzer SV 01" nation="GER">
          <CONTACT city="Mainz-Gonsenheim" country="DE" email="Guenter.Schmah@mainzersv01.de10" name="Schmah Günter" phone="06131-474854" state="RP" street="Max-Planck-Strasse 35c" zip="55124" />
          <ATHLETES>
            <ATHLETE birthdate="1938-01-01" firstname="Günter" gender="M" lastname="Schmah" nation="GER" license="12094" athleteid="6779">
              <ENTRIES>
                <ENTRY entrytime="00:01:35.00" eventid="1342" lane="5" heatid="8600" />
                <ENTRY entrytime="00:03:35.00" eventid="1304" lane="3" heatid="8583" />
                <ENTRY entrytime="00:00:40.00" eventid="1292" lane="6" heatid="8559" />
                <ENTRY entrytime="00:00:42.00" eventid="1284" lane="5" heatid="8546" />
                <ENTRY entrytime="00:01:36.00" eventid="1414" lane="3" heatid="8613" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1941-01-01" firstname="Franz" gender="M" lastname="Schlömer" nation="GER" license="12095" athleteid="6780">
              <ENTRIES>
                <ENTRY entrytime="00:01:42.00" eventid="1288" lane="4" heatid="8554" />
                <ENTRY entrytime="00:01:44.00" eventid="1296" lane="1" heatid="8565" />
                <ENTRY entrytime="00:03:38.00" eventid="1486" lane="3" heatid="8626" />
                <ENTRY entrytime="00:01:46.00" eventid="1414" lane="2" heatid="8613" />
                <ENTRY entrytime="00:00:42.00" eventid="1378" lane="3" heatid="8606" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCFG" name="SC Flipper Gossau" nation="SUI" region="ROS">
          <CONTACT city="Gossau" email="benedikt.rusch@helvetia.ch" fax="079 696 35 89" name="Rusch Benedikt" phone="058 280 43 65" street="Ilgenstrasse 7" zip="9200" />
          <ATHLETES>
            <ATHLETE birthdate="1954-01-01" firstname="Benedikt" gender="M" lastname="Rusch" nation="SUI" license="6282" athleteid="6792">
              <ENTRIES>
                <ENTRY entrytime="00:11:00.00" eventid="1196" lane="1" heatid="8590" />
                <ENTRY entrytime="00:00:34.00" eventid="1292" lane="4" heatid="8559" />
                <ENTRY entrytime="00:02:27.00" eventid="1107" lane="2" heatid="8540" />
                <ENTRY entrytime="00:05:16.00" eventid="1157" lane="3" heatid="8597" />
                <ENTRY entrytime="00:01:05.00" eventid="1450" lane="5" heatid="8623" />
                <ENTRY entrytime="00:02:55.00" eventid="1522" lane="2" heatid="8630" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SVE" name="Schwimmverein Emmen" nation="SUI" region="RZW">
          <ATHLETES>
            <ATHLETE birthdate="1962-10-12" firstname="Martin" gender="M" lastname="Grapentin" nation="SUI" license="25754" athleteid="6800">
              <ENTRIES>
                <ENTRY entrytime="00:02:40.00" eventid="1522" lane="3" heatid="8630" />
                <ENTRY entrytime="00:00:28.00" eventid="1300" lane="2" heatid="8580" />
                <ENTRY entrytime="00:00:30.00" eventid="1292" lane="5" heatid="8561" />
                <ENTRY entrytime="00:01:10.00" eventid="1342" lane="1" heatid="8601" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UET" name="SC Delphin Uetendorf" nation="SUI">
          <CONTACT city="Wattenwil" name="Berger Marianne" phone="033 356 24 38" street="Stafelalpstr.12" zip="3665" />
          <ATHLETES>
            <ATHLETE birthdate="1985-11-22" firstname="Nadja" gender="F" lastname="Bigler" nation="SUI" license="10084" athleteid="6807">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.80" eventid="1282" lane="4" heatid="8544" />
                <ENTRY entrytime="00:01:18.00" eventid="1294" lane="4" heatid="8564" />
                <ENTRY entrytime="00:01:24.50" eventid="1396" lane="3" heatid="8611" />
                <ENTRY entrytime="00:03:00.00" eventid="1302" lane="3" heatid="8582" />
                <ENTRY entrytime="00:05:00.00" eventid="1072" lane="2" heatid="8595" />
                <ENTRY entrytime="00:02:48.00" eventid="1504" lane="2" heatid="8629" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1989-10-06" firstname="Andrea" gender="F" lastname="Brechbühl" nation="SUI" license="15382" athleteid="6814">
              <ENTRIES>
                <ENTRY entrytime="00:02:50.00" eventid="1504" lane="5" heatid="8629" />
                <ENTRY entrytime="00:05:20.00" eventid="1072" lane="6" heatid="8595" />
                <ENTRY entrytime="00:01:14.00" eventid="1324" lane="2" heatid="8599" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-28" firstname="Yves" gender="M" lastname="Marclay" nation="SUI" license="3121" athleteid="6818">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.50" eventid="1288" lane="2" heatid="8556" />
                <ENTRY entrytime="00:00:32.00" eventid="1284" lane="1" heatid="8549" />
                <ENTRY entrytime="00:00:27.00" eventid="1300" lane="1" heatid="8581" />
                <ENTRY entrytime="00:01:09.50" eventid="1296" lane="6" heatid="8567" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCT" name="SC Thalwil" nation="SUI">
          <CONTACT city="Oberrieden" country="CH" email="heinzhaller@gmx.ch" name="Haller Heinz" street="Wiesengrundstr. 38" zip="8942" />
          <ATHLETES>
            <ATHLETE birthdate="1966-01-01" firstname="Robert" gender="M" lastname="Mundschin" nation="SUI" athleteid="6824">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.50" eventid="1292" lane="5" heatid="8560" />
                <ENTRY entrytime="00:00:28.50" eventid="1300" lane="3" heatid="8579" />
                <ENTRY entrytime="00:01:05.00" eventid="1450" lane="6" heatid="8623" />
                <ENTRY entrytime="00:02:27.00" eventid="1107" lane="4" heatid="8540" />
                <ENTRY entrytime="00:05:15.00" eventid="1157" lane="6" heatid="8598" />
                <ENTRY entrytime="00:00:38.00" eventid="1378" lane="1" heatid="8607" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Anja" gender="F" lastname="Gemperli" nation="SUI" athleteid="6887" />
            <ATHLETE birthdate="1959-01-01" firstname="Matthias" gender="M" lastname="Beusch" nation="SUI" athleteid="6888">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.50" eventid="1378" lane="6" heatid="8608" />
                <ENTRY entrytime="00:00:31.00" eventid="1292" lane="6" heatid="8561" />
                <ENTRY entrytime="00:00:29.00" eventid="1300" lane="3" heatid="8578" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Mauro" gender="M" lastname="Paulon" nation="SUI" athleteid="6889">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.00" eventid="1288" lane="2" heatid="8555" />
                <ENTRY entrytime="00:00:28.00" eventid="1300" lane="4" heatid="8580" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Fritz" gender="M" lastname="Keller" nation="SUI" athleteid="6890">
              <ENTRIES>
                <ENTRY entrytime="00:01:30.00" eventid="1450" lane="4" heatid="8621" />
                <ENTRY entrytime="00:01:37.00" eventid="1414" lane="4" heatid="8613" />
                <ENTRY entrytime="00:00:35.20" eventid="1300" lane="5" heatid="8576" />
                <ENTRY entrytime="00:00:42.50" eventid="1284" lane="6" heatid="8546" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Richard" gender="M" lastname="Niedermann" nation="SUI" athleteid="6891">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.82" eventid="1378" lane="3" heatid="8607" />
                <ENTRY entrytime="00:01:15.75" eventid="1288" lane="6" heatid="8556" />
                <ENTRY entrytime="00:00:28.65" eventid="1300" lane="2" heatid="8579" />
                <ENTRY entrytime="00:01:19.53" eventid="1296" lane="5" heatid="8566" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Manuel" gender="M" lastname="Strickler" nation="SUI" athleteid="6892">
              <ENTRIES>
                <ENTRY entrytime="00:01:18.00" eventid="1296" lane="2" heatid="8566" />
                <ENTRY entrytime="00:01:19.99" eventid="1414" lane="3" heatid="8614" />
                <ENTRY entrytime="00:01:21.00" eventid="1288" lane="5" heatid="8555" />
                <ENTRY entrytime="00:00:35.50" eventid="1284" lane="1" heatid="8548" />
                <ENTRY entrytime="00:00:36.00" eventid="1378" lane="5" heatid="8607" />
                <ENTRY entrytime="00:00:29.00" eventid="1300" lane="4" heatid="8578" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Arthur" gender="M" lastname="Rösler" nation="SUI" athleteid="6893">
              <ENTRIES>
                <ENTRY entrytime="00:06:10.00" eventid="1157" lane="3" heatid="8596" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Heinz" gender="M" lastname="Haller" nation="SUI" athleteid="6894">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.00" eventid="1284" lane="2" heatid="8547" />
                <ENTRY entrytime="00:00:32.50" eventid="1292" lane="4" heatid="8560" />
                <ENTRY entrytime="00:00:29.99" eventid="1300" lane="1" heatid="8578" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SV SS" name="Schwimmverein Sempachersee" nation="SUI">
          <CONTACT city="Willisau" country="CH" email="mcdiezi@bluemail.ch" name="Filli Martin" street="Höchhusmatt 19" zip="6030" />
          <ATHLETES>
            <ATHLETE birthdate="1939-01-01" firstname="Rene" gender="M" lastname="Diezi" nation="SUI" license="6098" athleteid="6826">
              <ENTRIES>
                <ENTRY entrytime="00:01:34.00" eventid="1296" lane="2" heatid="8565" />
                <ENTRY entrytime="00:01:38.00" eventid="1288" lane="3" heatid="8554" />
                <ENTRY entrytime="00:03:00.00" eventid="1107" lane="5" heatid="8539" />
                <ENTRY entrytime="00:04:00.00" eventid="1304" lane="2" heatid="8583" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1941-01-01" firstname="Maya-Claire" gender="F" lastname="Diezi" nation="SUI" license="445" athleteid="6827">
              <ENTRIES>
                <ENTRY entrytime="00:17:30.00" eventid="1177" lane="2" heatid="8587" />
                <ENTRY entrytime="00:04:50.00" eventid="1302" lane="5" heatid="8582" />
                <ENTRY entrytime="00:02:15.00" eventid="1294" lane="6" heatid="8563" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Simone" gender="F" lastname="Bürli" nation="SUI" athleteid="6926">
              <ENTRIES>
                <ENTRY entrytime="00:02:30.00" eventid="1054" lane="5" heatid="8537" />
                <ENTRY entrytime="00:10:30.00" eventid="1177" lane="4" heatid="8588" />
                <ENTRY entrytime="00:05:15.00" eventid="1072" lane="1" heatid="8595" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Martin" gender="M" lastname="Filli" nation="SUI" athleteid="6927">
              <ENTRIES>
                <ENTRY entrytime="00:01:25.00" eventid="1296" lane="3" heatid="8565" />
                <ENTRY entrytime="00:03:20.00" eventid="1522" lane="5" heatid="8630" />
                <ENTRY entrytime="00:11:30.00" eventid="1196" lane="4" heatid="8589" />
                <ENTRY entrytime="00:01:12.00" eventid="1450" lane="5" heatid="8622" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="Brigitte" gender="F" lastname="Herzog" nation="SUI" athleteid="6928">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.00" eventid="1298" lane="3" heatid="8571" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Bruno" gender="M" lastname="Moll" nation="SUI" athleteid="6929">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.00" eventid="1300" lane="4" heatid="8576" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="Andreas" gender="M" lastname="Moll" nation="SUI" athleteid="6930">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.00" eventid="1300" lane="6" heatid="8576" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-16" firstname="Bertrand" gender="M" lastname="Grob" nation="SUI" athleteid="7878">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.50" eventid="1292" lane="3" heatid="8560" />
                <ENTRY entrytime="00:00:36.00" eventid="1284" lane="6" heatid="8548" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Heidi" gender="F" lastname="Arnold" nation="SUI" athleteid="8710" />
            <ATHLETE birthdate="1969-12-25" firstname="Andreas" gender="M" lastname="Murer" nation="SUI" athleteid="8711" />
            <ATHLETE firstname="Martin" gender="M" lastname="Grapentin" nation="SUI" athleteid="10220" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1175" lane="6" heatid="8585">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6928" number="1" />
                    <RELAYPOSITION athleteid="7878" number="2" />
                    <RELAYPOSITION athleteid="6926" number="3" />
                    <RELAYPOSITION athleteid="6927" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="NT" eventid="1540" lane="1" heatid="8633">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6800" number="1" />
                    <RELAYPOSITION athleteid="6926" number="2" />
                    <RELAYPOSITION athleteid="8710" number="3" />
                    <RELAYPOSITION athleteid="6927" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1175" lane="1" heatid="8585">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6827" number="1" />
                    <RELAYPOSITION athleteid="8710" number="2" />
                    <RELAYPOSITION athleteid="6826" number="3" />
                    <RELAYPOSITION athleteid="8711" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="RFN" name="Red Fish Neuchatel" nation="SUI" region="RSR">
          <ATHLETES>
            <ATHLETE birthdate="1966-07-21" firstname="Claudia" gender="F" lastname="Lautenbacher" nation="SUI" athleteid="6836">
              <ENTRIES>
                <ENTRY entrytime="00:02:48.00" eventid="1504" lane="4" heatid="8629" />
                <ENTRY entrytime="00:01:25.00" eventid="1396" lane="4" heatid="8611" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1966-09-17" firstname="Philippe" gender="M" lastname="Allegrini" nation="SUI" license="2383" athleteid="7283">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1196" lane="3" heatid="9736" />
                <ENTRY entrytime="NT" eventid="7347" lane="4" heatid="8592" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LN" name="Lausanne Natation" nation="SUI" region="RSR">
          <CONTACT city="Lausanne" email="cedric.cattaneo@gmail.com" fax="0216165160" name="Cattaneo Cédric" phone="0216165159" state="VD" street="Av. du Servan 32" zip="1006" />
          <ATHLETES>
            <ATHLETE birthdate="1984-07-04" firstname="Sébastien" gender="M" lastname="Boutinard Rouelle" nation="SUI" athleteid="6840">
              <ENTRIES>
                <ENTRY entrytime="00:00:43.00" eventid="1378" lane="2" heatid="8606" />
                <ENTRY entrytime="00:01:04.00" eventid="1450" lane="6" heatid="8624" />
                <ENTRY entrytime="00:00:28.50" eventid="1300" lane="1" heatid="8580" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1972-05-25" firstname="Rainer" gender="M" lastname="Buchholz" nation="GER" athleteid="6844">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.50" eventid="1300" lane="2" heatid="8581" />
                <ENTRY entrytime="00:01:04.00" eventid="1288" lane="4" heatid="8556" />
                <ENTRY entrytime="00:00:57.50" eventid="1450" status="WDR" />
                <ENTRY entrytime="00:00:29.50" eventid="1378" status="WDR" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-26" firstname="Cédric" gender="M" lastname="Cattaneo" nation="SUI" athleteid="6849">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.90" eventid="1450" status="WDR" />
                <ENTRY entrytime="00:01:19.50" eventid="1414" status="WDR" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-05" firstname="Eavan" gender="F" lastname="Dorcey" nation="IRL" athleteid="6854" />
            <ATHLETE birthdate="1989-05-10" firstname="Agustin" gender="M" lastname="Gutierrez" nation="SUI" athleteid="6858">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="1450" lane="4" heatid="8623" />
                <ENTRY entrytime="00:00:36.00" eventid="1284" lane="3" heatid="8547" />
                <ENTRY entrytime="00:01:20.00" eventid="1414" lane="2" heatid="8614" />
                <ENTRY entrytime="00:00:28.50" eventid="1300" lane="4" heatid="8579" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-21" firstname="Osamu" gender="M" lastname="Moser" nation="SUI" athleteid="6863">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.00" eventid="1414" lane="1" heatid="8615" />
                <ENTRY entrytime="00:01:07.00" eventid="1296" lane="5" heatid="8567" />
                <ENTRY entrytime="00:00:32.00" eventid="1284" lane="5" heatid="8549" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-21" firstname="Nicole" gender="F" lastname="Solenthaler" nation="SUI" athleteid="6867">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.50" eventid="1360" lane="4" heatid="8604" />
                <ENTRY entrytime="00:01:24.00" eventid="1286" lane="4" heatid="8552" />
                <ENTRY entrytime="00:01:16.00" eventid="1432" lane="4" heatid="8618" />
                <ENTRY entrytime="00:01:24.00" eventid="1294" lane="1" heatid="8564" />
                <ENTRY entrytime="00:00:33.00" eventid="1298" lane="1" heatid="8573" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-16" firstname="David" gender="M" lastname="Tron" nation="LUX" athleteid="6873">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.50" eventid="1378" lane="1" heatid="8608" />
                <ENTRY entrytime="00:01:08.00" eventid="1296" lane="1" heatid="8567" />
                <ENTRY entrytime="00:00:59.50" eventid="1450" lane="2" heatid="8624" />
                <ENTRY entrytime="00:00:27.00" eventid="1300" lane="6" heatid="8581" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1990-04-10" firstname="Moira" gender="F" lastname="Wacker" nation="SUI" athleteid="6878">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.00" eventid="1298" lane="4" heatid="8572" />
                <ENTRY entrytime="00:01:32.00" eventid="1396" lane="5" heatid="8611" />
                <ENTRY entrytime="00:00:43.00" eventid="1282" lane="2" heatid="8544" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:30.00" eventid="1175" lane="5" heatid="8585">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6867" number="1" />
                    <RELAYPOSITION athleteid="6878" number="2" />
                    <RELAYPOSITION athleteid="6844" number="3" />
                    <RELAYPOSITION athleteid="6840" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:02:10.00" eventid="1540" lane="2" heatid="8633">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6858" number="1" />
                    <RELAYPOSITION athleteid="6867" number="2" />
                    <RELAYPOSITION athleteid="6878" number="3" />
                    <RELAYPOSITION athleteid="6873" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AARE" name="Schwimmclub Aarefisch" nation="SUI">
          <CONTACT city="Aarau" email="samuel..nikles@bluewin.ch" street="Weihermattstr. 74/76" zip="5000" />
          <ATHLETES>
            <ATHLETE birthdate="1984-02-14" firstname="Samuel" gender="M" lastname="Niklès" nation="SUI" athleteid="6885">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.45" eventid="1300" lane="3" heatid="8575" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-04" firstname="Alfonso" gender="M" lastname="Die" nation="SUI" athleteid="8635">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1300" lane="1" heatid="8574" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TMJPN" name="Tousuikai Masters" nation="JPN">
          <CONTACT city="Brugg" country="CH" email="Yohei.Sato@psi.ch" name="Yohei Sato" street="Sommerhaldenstrasse 1a" zip="5200" />
          <ATHLETES>
            <ATHLETE birthdate="1972-09-14" firstname="Yohei" gender="M" lastname="Sato" nation="JPN" license="13-110" athleteid="6942" externalid="720914-2">
              <ENTRIES>
                <ENTRY entrytime="00:02:27.00" eventid="1522" lane="2" heatid="8631" />
                <ENTRY entrytime="00:01:20.00" eventid="1414" lane="4" heatid="8614" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SVB" name="Schwimmverein beider Basel" nation="SUI" region="RZW">
          <CONTACT city="Therwil" email="mtolusso@hotmail.com" name="Tolusso Markus" phone="061 721 00 52" street="Teichstrasse 47" zip="4106" />
          <ATHLETES>
            <ATHLETE birthdate="1976-04-23" firstname="Peter" gender="M" lastname="Bezak" nation="SUI" license="279" athleteid="6946">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="1450" lane="2" heatid="8623" />
                <ENTRY entrytime="00:00:31.00" eventid="1292" lane="1" heatid="8561" />
                <ENTRY entrytime="00:05:05.00" eventid="1157" lane="5" heatid="8598" />
                <ENTRY entrytime="00:00:29.50" eventid="1300" lane="2" heatid="8578" />
                <ENTRY entrytime="00:00:38.00" eventid="1284" lane="5" heatid="8547" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1963-09-17" firstname="Roger" gender="M" lastname="Birrer" nation="SUI" athleteid="6952">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.00" eventid="1378" lane="3" heatid="8608" />
                <ENTRY entrytime="00:01:01.50" eventid="1342" lane="4" heatid="8601" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-02" firstname="Stefan" gender="M" lastname="Brand" nation="SUI" license="8010" athleteid="6958">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.50" eventid="1292" lane="3" heatid="8561" />
                <ENTRY entrytime="00:00:53.00" eventid="1450" lane="3" heatid="8624" />
                <ENTRY entrytime="00:00:59.90" eventid="1342" lane="3" heatid="8601" />
                <ENTRY entrytime="00:00:24.50" eventid="1300" lane="4" heatid="8581" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Heidi" gender="F" lastname="Clark" nation="SUI" athleteid="6963">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.00" eventid="1298" lane="6" heatid="8573" />
                <ENTRY entrytime="00:01:10.00" eventid="1432" lane="1" heatid="8619" />
                <ENTRY entrytime="00:05:45.00" eventid="1072" lane="4" heatid="8594" />
                <ENTRY entrytime="00:02:45.00" eventid="1054" lane="4" heatid="8536" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-03" firstname="Margarethe" gender="F" lastname="Denk" nation="GER" license="18490" athleteid="6966">
              <ENTRIES>
                <ENTRY entrytime="00:01:21.00" eventid="1324" lane="5" heatid="8599" />
                <ENTRY entrytime="00:12:07.00" eventid="1177" lane="5" heatid="8588" />
                <ENTRY entrytime="00:01:22.00" eventid="1294" lane="5" heatid="8564" />
                <ENTRY entrytime="00:00:35.00" eventid="1290" lane="4" heatid="8557" />
                <ENTRY entrytime="00:03:15.00" eventid="1504" lane="2" heatid="8628" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1946-09-26" firstname="Kurt" gender="M" lastname="Frei" nation="SUI" license="4468" athleteid="6972">
              <ENTRIES>
                <ENTRY entrytime="00:02:50.00" eventid="1486" lane="5" heatid="8627" />
                <ENTRY entrytime="00:00:36.00" eventid="1378" lane="2" heatid="8607" />
                <ENTRY entrytime="00:01:15.00" eventid="1288" lane="1" heatid="8556" />
                <ENTRY entrytime="00:05:40.00" eventid="1157" lane="2" heatid="8597" />
                <ENTRY entrytime="00:11:30.00" eventid="1196" lane="3" heatid="8589" />
                <ENTRY entrytime="00:00:31.00" eventid="1300" lane="5" heatid="8577" />
                <ENTRY entrytime="00:02:30.00" eventid="1107" lane="1" heatid="8540" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-10" firstname="Irene" gender="F" lastname="Nestor" nation="SUI" license="607" athleteid="6980">
              <ENTRIES>
                <ENTRY entrytime="00:01:32.00" eventid="1286" lane="3" heatid="8551" />
                <ENTRY entrytime="00:02:56.00" eventid="1054" lane="5" heatid="8536" />
                <ENTRY entrytime="00:01:35.00" eventid="1294" lane="4" heatid="8563" />
                <ENTRY entrytime="00:03:14.00" eventid="1468" lane="4" heatid="8625" />
                <ENTRY entrytime="00:12:25.00" eventid="1177" lane="3" heatid="8587" />
                <ENTRY entrytime="00:06:10.00" eventid="1072" lane="1" heatid="8594" />
                <ENTRY entrytime="00:00:45.00" eventid="1360" lane="6" heatid="8604" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1955-12-14" firstname="Ferdy" gender="M" lastname="Polasek" nation="SUI" license="16664" athleteid="6988">
              <ENTRIES>
                <ENTRY entrytime="00:05:15.00" eventid="1157" lane="1" heatid="8598" />
                <ENTRY entrytime="00:02:25.00" eventid="1107" lane="3" heatid="8540" />
                <ENTRY entrytime="00:00:40.00" eventid="1284" lane="3" heatid="8546" />
                <ENTRY entrytime="00:11:00.00" eventid="1196" lane="6" heatid="8590" />
                <ENTRY entrytime="00:01:06.00" eventid="1450" lane="3" heatid="8622" />
                <ENTRY entrytime="00:00:29.90" eventid="1300" lane="5" heatid="8578" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1949-05-30" firstname="Mireille" gender="F" lastname="Richter" nation="SUI" license="5930" athleteid="6995">
              <ENTRIES>
                <ENTRY entrytime="00:01:57.50" eventid="1396" lane="2" heatid="8610" />
                <ENTRY entrytime="00:03:09.00" eventid="1054" lane="3" heatid="8535" />
                <ENTRY entrytime="00:03:59.00" eventid="1302" lane="4" heatid="8582" />
                <ENTRY entrytime="NT" eventid="1177" lane="5" heatid="8587" />
                <ENTRY entrytime="00:24:17.00" eventid="7347" lane="3" heatid="8592" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-15" firstname="Regula" gender="F" lastname="Steiger" nation="SUI" license="514" athleteid="7000">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.50" eventid="1298" lane="4" heatid="8573" />
                <ENTRY entrytime="00:01:26.00" eventid="1396" lane="2" heatid="8611" />
                <ENTRY entrytime="00:00:38.80" eventid="1282" lane="3" heatid="8544" />
                <ENTRY entrytime="00:01:08.00" eventid="1432" status="DNS" lane="5" heatid="8619" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1958-08-10" firstname="Markus" gender="M" lastname="Tolusso" nation="SUI" athleteid="7005">
              <ENTRIES>
                <ENTRY entrytime="00:01:30.00" eventid="1288" lane="6" heatid="8555" />
                <ENTRY entrytime="00:01:30.00" eventid="1296" lane="4" heatid="8565" />
                <ENTRY entrytime="00:00:34.00" eventid="1292" lane="6" heatid="8560" />
                <ENTRY entrytime="00:12:00.00" eventid="1196" lane="2" heatid="8589" />
                <ENTRY entrytime="00:00:32.50" eventid="1300" lane="3" heatid="8576" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.00" eventid="1540" lane="4" heatid="8633">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6946" number="1">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="6963" number="2">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="6988" number="3">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="6966" number="4">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:02:07.80" eventid="1175" lane="4" heatid="8585">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6972" number="1">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="7000" number="2">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="6958" number="3">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="6963" number="4">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SRM" name="SK Region Murten" nation="SUI" region="RSR">
          <CONTACT city="Murten" email="keiju@bluewin.ch" name="Herzig Heidi" street="Prehlstr. 35" zip="3280" />
          <ATHLETES>
            <ATHLETE birthdate="1966-04-17" firstname="Alexis" gender="M" lastname="Bögli" nation="SUI" license="12118" athleteid="7081">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.50" eventid="1284" lane="6" heatid="8549" />
                <ENTRY entrytime="00:01:14.00" eventid="1414" lane="5" heatid="8615" />
                <ENTRY entrytime="00:04:55.00" eventid="1157" lane="2" heatid="8598" />
                <ENTRY entrytime="00:00:27.90" eventid="1300" lane="3" heatid="8580" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1960-07-30" firstname="Anita" gender="F" lastname="Zingg" nation="SUI" license="4769" athleteid="7086">
              <ENTRIES>
                <ENTRY entrytime="00:01:22.00" eventid="1286" lane="3" heatid="8552" />
                <ENTRY entrytime="00:02:38.00" eventid="1054" lane="1" heatid="8537" />
                <ENTRY entrytime="00:05:30.00" eventid="1072" status="WDR" />
                <ENTRY entrytime="00:01:10.00" eventid="1432" status="WDR" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WITT" name="Schwimm-Club Wittenbach" nation="SUI" region="ROS">
          <CONTACT city="St.Gallen" email="gabschneider@gmx.net" name="Schneider Gabriel" street="Lukasstr.5" zip="9008" />
          <ATHLETES>
            <ATHLETE birthdate="1972-11-11" firstname="Matthias" gender="M" lastname="Baumberger" nation="SUI" license="23131" athleteid="7092">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="1450" status="WDR" />
                <ENTRY entrytime="00:05:45.00" eventid="1157" status="WDR" />
                <ENTRY entrytime="00:00:31.13" eventid="1300" status="WDR" />
                <ENTRY entrytime="00:02:34.00" eventid="1107" status="WDR" />
                <ENTRY entrytime="00:00:37.27" eventid="1292" status="WDR" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PLAN" name="CN Plan-les-Ouates" nation="SUI" region="RSR">
          <CONTACT city="Châtelaine" email="rascha54@yahoo.fr" name="Schallon Ralph" phone="022 796 79 83" street="av. de Crozet 12" street2="Directeur technique" zip="1219" />
          <ATHLETES>
            <ATHLETE birthdate="1953-06-12" firstname="Alexandre" gender="M" lastname="Barrena" nation="SUI" license="13184" athleteid="7099" />
            <ATHLETE birthdate="1965-07-13" firstname="Murielle" gender="F" lastname="Caillet Dayer" nation="SUI" license="1035" athleteid="7102">
              <ENTRIES>
                <ENTRY entrytime="00:01:32.28" eventid="1286" lane="4" heatid="8551">
                  <MEETINFO city="Plan-les-Ouates" course="SCM" date="2009-03-14" name="Masters Meet PLO" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:03:10.00" eventid="1468" lane="3" heatid="8625" />
                <ENTRY entrytime="00:00:40.90" eventid="1360" lane="5" heatid="8604" />
                <ENTRY entrytime="00:00:37.00" eventid="1298" lane="6" heatid="8572" />
                <ENTRY entrytime="00:01:35.00" eventid="1294" lane="5" heatid="8563" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1963-12-23" firstname="Patricia" gender="F" lastname="Kamm" nation="SUI" license="24901" athleteid="7108">
              <ENTRIES>
                <ENTRY entrytime="00:12:46.27" eventid="1177" lane="4" heatid="8587">
                  <MEETINFO city="Oerlikon" course="LCM" date="2009-08-23" name="2. Zurich International Masters Championships" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:06:11.42" eventid="1072" lane="3" heatid="8593">
                  <MEETINFO city="Oerlikon" course="LCM" date="2009-08-22" name="2. Zurich International Masters Championships" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.40" eventid="1432" lane="5" heatid="8618">
                  <MEETINFO city="Ferney-Voltaire" course="SCM" date="2009-06-13" name="Coupe de l&apos;Ain des Maîtres" nation="FRA" />
                </ENTRY>
                <ENTRY entrytime="00:01:26.33" eventid="1286" lane="2" heatid="8552">
                  <MEETINFO city="Ferney-Voltaire" course="SCM" date="2009-06-13" name="Coupe de l&apos;Ain des Maîtres" nation="FRA" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1965-07-21" firstname="Nathalie" gender="F" lastname="Landenbergue" nation="SUI" license="1736" athleteid="7113">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.85" eventid="1298" lane="2" heatid="8572">
                  <MEETINFO city="Plan-les-Ouates" course="SCM" date="2008-10-11" name="Championnat interne 2008" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.02" eventid="1282" lane="5" heatid="8544">
                  <MEETINFO city="Plan-les-Ouates" course="SCM" date="2008-10-11" name="Championnat interne 2008" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.14" eventid="1432" lane="2" heatid="8618">
                  <MEETINFO city="Belfort" course="SCM" date="2008-11-30" name="2e Challenge 4-nages des Maîtres" nation="FRA" />
                </ENTRY>
                <ENTRY entrytime="00:01:36.62" eventid="1396" lane="1" heatid="8611">
                  <MEETINFO city="Plan-les-Ouates" course="SCM" date="2009-03-14" name="Masters Meet PLO" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.58" eventid="1294" lane="6" heatid="8564">
                  <MEETINFO city="Belfort" course="SCM" date="2008-11-30" name="2e Challenge 4-nages des Maîtres" nation="FRA" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1969-08-15" firstname="Xavier" gender="M" lastname="Louis" nation="SUI" license="23189" athleteid="7119">
              <ENTRIES>
                <ENTRY entrytime="00:01:18.96" eventid="1288" lane="4" heatid="8555">
                  <MEETINFO city="Genève" course="SCM" date="2009-01-24" name="2ème Meeting Inter-Clubs NSG saison 2008-2009" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.00" eventid="1486" lane="1" heatid="8627" />
                <ENTRY entrytime="00:00:34.88" eventid="1378" lane="4" heatid="8607">
                  <MEETINFO city="Le Fayet" course="SCM" date="2009-05-16" name="Marathons du Mont-Blanc" nation="FRA" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.90" eventid="1300" lane="6" heatid="8579">
                  <MEETINFO city="Plan-les-Ouates" course="SCM" date="2009-03-14" name="Masters Meet PLO" nation="SUI" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-03" firstname="Antoine" gender="M" lastname="Mayerat" nation="SUI" license="26076" athleteid="7124">
              <ENTRIES>
                <ENTRY entrytime="00:02:40.00" eventid="1522" lane="6" heatid="8631">
                  <MEETINFO city="Plan-les-Ouates" course="SCM" date="2009-06-18" name="Test interne" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.81" eventid="1342" lane="6" heatid="8601">
                  <MEETINFO city="Ferney-Voltaire" course="SCM" date="2009-06-13" name="Coupe de l&apos;Ain des Maîtres" nation="FRA" />
                </ENTRY>
                <ENTRY entrytime="00:09:45.00" eventid="1196" lane="4" heatid="8590" />
                <ENTRY entrytime="00:01:03.50" eventid="1450" lane="1" heatid="8624">
                  <MEETINFO city="Ferney-Voltaire" course="SCM" date="2009-06-13" name="Coupe de l&apos;Ain des Maîtres" nation="FRA" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.00" eventid="1107" lane="2" heatid="8541" />
                <ENTRY entrytime="00:00:32.82" eventid="1292" lane="2" heatid="8560">
                  <MEETINFO city="Annemasse" course="SCM" date="2009-04-04" name="Meeting Masters" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.89" eventid="1300" lane="1" heatid="8579">
                  <MEETINFO city="Ferney-Voltaire" course="SCM" date="2009-06-13" name="Coupe de l&apos;Ain des Maîtres" nation="FRA" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1954-07-02" firstname="Ralph" gender="M" lastname="Schallon" nation="SUI" license="3101" athleteid="7132">
              <ENTRIES>
                <ENTRY entrytime="00:02:45.95" eventid="1304" lane="2" heatid="8584">
                  <MEETINFO city="Belfort" course="SCM" date="2008-11-30" name="2e Challenge 4-nages des Maîtres" nation="FRA" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.76" eventid="1414" lane="6" heatid="8615">
                  <MEETINFO city="Plan-les-Ouates" course="SCM" date="2009-03-26" name="Test interne brasse" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.81" eventid="1284" lane="2" heatid="8548">
                  <MEETINFO city="Plan-les-Ouates" course="SCM" date="2009-03-14" name="Masters Meet PLO" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.00" eventid="1522" lane="4" heatid="8630" />
                <ENTRY entrytime="00:01:13.20" eventid="1296" status="WDR">
                  <MEETINFO city="Plan-les-Ouates" course="SCM" date="2009-03-14" name="Masters Meet PLO" nation="SUI" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:02:17.51" eventid="1540" lane="5" heatid="8633">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7119" number="1">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="7108" number="2">
                      <MEETINFO city="Ferney-Voltaire" course="SCM" date="2009-06-13" name="Coupe de l&apos;Ain des Maîtres" nation="FRA" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="7113" number="3">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="7124" number="4">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:02:27.20" eventid="1175" lane="2" heatid="8585">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7102" number="1">
                      <MEETINFO city="Le Fayet" course="SCM" date="1909-05-16" name="Marathons du Mont-Blanc" nation="FRA" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="7132" number="2">
                      <MEETINFO city="Plan-les-Ouates" course="SCM" date="1908-10-11" name="Championnat interne 2008" nation="SUI" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="7119" number="3">
                      <MEETINFO city="Annemasse" course="SCM" date="1909-04-04" name="Meeting Masters" />
                    </RELAYPOSITION>
                    <RELAYPOSITION athleteid="7113" number="4">
                      <MEETINFO course="SCM" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AVU" name="Avully Natation" nation="SUI" region="RSR">
          <CONTACT city="Sézegnin" name="Gaspoz Olivier" phone="022 756 20 94" street="33 rte du Creux-du-Loup" zip="1285" />
          <ATHLETES>
            <ATHLETE birthdate="1973-08-24" firstname="Laurent" gender="M" lastname="Thévenaz" nation="SUI" license="17578" athleteid="7139">
              <ENTRIES>
                <ENTRY entrytime="00:02:35.00" eventid="1486" lane="2" heatid="8627" />
                <ENTRY entrytime="00:04:55.00" eventid="1157" lane="4" heatid="8598" />
                <ENTRY entrytime="00:10:30.00" eventid="1196" lane="5" heatid="8590" />
                <ENTRY entrytime="00:02:15.00" eventid="1107" lane="5" heatid="8541" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BREM" name="SC Region Bremgarten" nation="SUI" region="RZO">
          <CONTACT city="Bremgarten 2" email="info@scrb.ch" internet="www.scrb.ch" name="Andy Kempter" street2="Postfach 2123" zip="5620" />
          <ATHLETES>
            <ATHLETE birthdate="1957-07-30" firstname="Brigitte" gender="F" lastname="Christen" nation="SUI" license="22603" athleteid="7147">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.50" eventid="1298" lane="1" heatid="8571" />
                <ENTRY entrytime="00:03:52.00" eventid="1054" lane="4" heatid="8535" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Matthias" gender="M" lastname="Fehlmann" nation="SUI" athleteid="7150">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.49" eventid="1284" lane="6" heatid="8547">
                  <MEETINFO city="78050 Villingen-Schwenningen" course="SCM" date="2009-04-04" name="36. Internationale Masters-Meeting des Schwimm-Club-Villingen von 1950 e.V." nation="GER" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="1107" lane="2" heatid="8538" />
                <ENTRY entrytime="00:00:32.22" eventid="1300" status="WDR" lane="6" heatid="8577">
                  <MEETINFO city="78050 Villingen-Schwenningen" course="SCM" date="1909-04-04" name="36. Internationale Masters-Meeting des Schwimm-Club-Villingen von 1950 e.V." nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:03:25.00" eventid="1304" status="WDR" lane="6" heatid="8584" />
                <ENTRY entrytime="00:01:28.25" eventid="1414" status="WDR">
                  <MEETINFO city="78050 Villingen-Schwenningen" course="SCM" date="1909-04-04" name="36. Internationale Masters-Meeting des Schwimm-Club-Villingen von 1950 e.V." nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.53" eventid="1450" status="WDR">
                  <MEETINFO city="78050 Villingen-Schwenningen" course="SCM" date="1909-04-04" name="36. Internationale Masters-Meeting des Schwimm-Club-Villingen von 1950 e.V." nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1958-12-06" firstname="Andy" gender="M" lastname="Kempter" nation="SUI" athleteid="7157">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.56" eventid="1378" lane="4" heatid="8606" />
                <ENTRY entrytime="00:01:22.36" eventid="1450" lane="3" heatid="8621" />
                <ENTRY entrytime="00:00:47.75" eventid="1292" lane="4" heatid="8558" />
                <ENTRY entrytime="00:00:34.29" eventid="1300" lane="2" heatid="8576" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1960-08-09" firstname="Melanie" gender="F" lastname="Lins" nation="SUI" athleteid="7162">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.00" eventid="1282" lane="4" heatid="8543" />
                <ENTRY entrytime="00:00:41.00" eventid="1298" lane="5" heatid="8571" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1956-02-21" firstname="Ruth" gender="F" lastname="Stierli" nation="SUI" license="22083" athleteid="7165">
              <ENTRIES>
                <ENTRY entrytime="00:04:10.00" eventid="1302" lane="2" heatid="8582" />
                <ENTRY entrytime="00:00:48.74" eventid="1282" lane="3" heatid="8543">
                  <MEETINFO city="78050 Villingen-Schwenningen" course="SCM" date="2009-04-04" name="36. Internationale Masters-Meeting des Schwimm-Club-Villingen von 1950 e.V." nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Paul" gender="M" lastname="Spadt" nation="SUI" athleteid="7872">
              <ENTRIES>
                <ENTRY entrytime="00:02:27.00" eventid="1522" lane="5" heatid="8631" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BUEL" name="Schwimmclub Bülach" nation="SUI" region="RZO">
          <CONTACT city="Windlach" email="tibi.kiss@bluewin.ch" name="Kiss Tibor" phone="01/862 6001" street="Raaterstr. 20" zip="8175" />
          <ATHLETES>
            <ATHLETE birthdate="1983-03-01" firstname="Andrea" gender="F" lastname="Bächli" nation="SUI" license="10378" athleteid="7169">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.94" eventid="1294" lane="2" heatid="8564">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:10:18.96" eventid="1177" lane="3" heatid="8588">
                  <MEETINFO city="Oerlikon" course="LCM" date="2009-08-23" name="2. Zurich International Masters Championships" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.58" eventid="1432" lane="4" heatid="8619">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.38" eventid="1054" lane="4" heatid="8537">
                  <MEETINFO city="Hallenbad Biel-Bienne" course="SCM" date="1909-05-02" name="Bieler Nachwuchs-Wettkämpfe 2009" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:04:57.70" eventid="1072" lane="4" heatid="8595">
                  <MEETINFO city="Hallenbad Biel-Bienne" course="SCM" date="2009-05-03" name="Bieler Nachwuchs-Wettkämpfe 2009" nation="SUI" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-10" firstname="Patrice" gender="M" lastname="Pellaton" nation="SUI" license="1722" athleteid="7175">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.07" eventid="1107" lane="4" heatid="8541">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.24" eventid="1300" lane="3" heatid="8581">
                  <MEETINFO city="Lausanne" course="SCM" date="2008-11-28" name="FSN: Kurzbahn - Schweizermeisterschaft" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.80" eventid="1292" lane="2" heatid="8561">
                  <MEETINFO city="Lausanne" course="SCM" date="2008-11-30" name="FSN: Kurzbahn - Schweizermeisterschaft" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.00" eventid="1450" lane="4" heatid="8624">
                  <MEETINFO city="Lausanne" course="SCM" date="2008-11-30" name="FSN: Kurzbahn - Schweizermeisterschaft" nation="SUI" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.25" eventid="1342" lane="2" heatid="8601">
                  <MEETINFO city="Hallenbad Biel-Bienne" course="SCM" date="2009-01-31" name="Meeting Intervilles 2009" nation="SUI" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1965-10-14" firstname="Alfredo" gender="M" lastname="Prencipe" nation="GER" athleteid="7181">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.59" eventid="1450" lane="3" heatid="8623" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="HSV" name="HSV Medizin Magdeburg" nation="GER">
          <CONTACT city="Magdeburg" email="klesinski@email.de" name="Gerald Schmidt" street="Hannoversche Str. 7d" zip="39110" />
          <ATHLETES>
            <ATHLETE birthdate="1976-09-22" firstname="René" gender="M" lastname="Klesinski" nation="GER" license="074167" athleteid="7184">
              <ENTRIES>
                <ENTRY entrytime="00:02:19.21" eventid="1107" lane="1" heatid="8541" />
                <ENTRY entrytime="00:00:34.21" eventid="1292" lane="2" heatid="8559" />
                <ENTRY entrytime="00:01:15.99" eventid="1288" lane="3" heatid="8555" />
                <ENTRY entrytime="00:00:28.87" eventid="1300" lane="5" heatid="8579" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AMT" name="Aquatic Masters Team" nation="SUI">
          <CONTACT city="Bollingen" email="cristian58@bluewin.ch" name="Cristian Rentsch" street="Dorfstrasse 55" zip="8715" />
          <ATHLETES>
            <ATHLETE birthdate="1969-01-01" firstname="Basil" gender="M" lastname="Düby" nation="SUI" athleteid="7190">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="1342" lane="5" heatid="8601" />
                <ENTRY entrytime="00:02:35.00" eventid="1522" lane="1" heatid="8631" />
                <ENTRY entrytime="00:01:05.00" eventid="1450" lane="1" heatid="8623" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Toni" gender="M" lastname="Pavicic-Donkic" nation="SUI" license="10982" athleteid="7191">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.12" eventid="1107" lane="3" heatid="8541" />
                <ENTRY entrytime="00:04:14.92" eventid="1157" lane="3" heatid="8598" />
                <ENTRY entrytime="00:02:24.10" eventid="1522" lane="4" heatid="8631" />
                <ENTRY entrytime="00:08:59.70" eventid="1196" status="DNS" lane="3" heatid="8590" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Christian" gender="M" lastname="Rentsch" nation="SUI" license="843" athleteid="7192">
              <ENTRIES>
                <ENTRY entrytime="00:02:43.00" eventid="1304" lane="4" heatid="8584" />
                <ENTRY entrytime="00:02:30.00" eventid="1486" lane="3" heatid="8627" />
                <ENTRY entrytime="00:00:33.00" eventid="1284" lane="4" heatid="8548" />
                <ENTRY entrytime="00:05:25.00" eventid="1157" status="DNS" lane="4" heatid="8597" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Sonja" gender="F" lastname="Gwerder" nation="SUI" license="13520" athleteid="7193">
              <ENTRIES>
                <ENTRY entrytime="00:02:40.00" eventid="1504" lane="3" heatid="8629" />
                <ENTRY entrytime="00:01:13.00" eventid="1294" lane="3" heatid="8564" />
                <ENTRY entrytime="00:01:11.00" eventid="1324" lane="4" heatid="8599" />
                <ENTRY entrytime="00:00:34.00" eventid="1360" lane="3" heatid="8604" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Alicia" gender="F" lastname="Irvin" nation="SUI" license="13815" athleteid="7194">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.00" eventid="1298" lane="3" heatid="8573" />
                <ENTRY entrytime="00:02:50.00" eventid="1054" lane="2" heatid="8536" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Evgenia" gender="F" lastname="Bedenig" nation="SUI" athleteid="7195">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.00" eventid="1290" lane="3" heatid="8557" />
                <ENTRY entrytime="00:01:10.00" eventid="1324" lane="3" heatid="8599" />
                <ENTRY entrytime="00:01:05.00" eventid="1432" lane="3" heatid="8619" />
                <ENTRY entrytime="00:02:20.00" eventid="1054" lane="3" heatid="8537" />
                <ENTRY entrytime="00:04:40.00" eventid="1072" lane="3" heatid="8595" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.00" eventid="1175" lane="3" heatid="8585">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7192" number="1" />
                    <RELAYPOSITION athleteid="7191" number="2" />
                    <RELAYPOSITION athleteid="7193" number="3" />
                    <RELAYPOSITION athleteid="7194" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <ENTRIES>
                <ENTRY entrytime="00:01:52.00" eventid="1540" lane="3" heatid="8633">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7190" number="1" />
                    <RELAYPOSITION athleteid="7191" number="2" />
                    <RELAYPOSITION athleteid="7193" number="3" />
                    <RELAYPOSITION athleteid="7195" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TSV" name="TSV 1862 Erding" nation="GER">
          <CONTACT email="delphine.erding@t-online.de" name="Petra Teichert" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Hans Georg" gender="M" lastname="Fiedeldeij" nation="GER" license="154290" athleteid="7201">
              <ENTRIES>
                <ENTRY entrytime="00:10:24.42" eventid="1196" lane="2" heatid="8590" />
                <ENTRY entrytime="00:00:28.16" eventid="1300" lane="5" heatid="8580" />
                <ENTRY entrytime="00:02:19.60" eventid="1107" lane="6" heatid="8541" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCW" name="SC Winterthur" nation="SUI">
          <CONTACT email="mueller.peter@bluewin.ch" name="Peter Müller" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Markus" gender="M" lastname="Enz" nation="SUI" license="715" athleteid="7203">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.00" eventid="1296" lane="1" heatid="8566" />
                <ENTRY entrytime="00:02:30.00" eventid="1107" lane="6" heatid="8540" />
                <ENTRY entrytime="00:00:35.00" eventid="1292" lane="5" heatid="8559" />
                <ENTRY entrytime="00:00:30.50" eventid="1300" lane="6" heatid="8578" />
                <ENTRY entrytime="00:00:39.00" eventid="1284" lane="1" heatid="8547" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Marcel" gender="M" lastname="Schwarz" nation="SUI" license="8657" athleteid="7204">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.00" eventid="1284" lane="3" heatid="8548" />
                <ENTRY entrytime="00:00:28.50" eventid="1300" lane="6" heatid="8580" />
                <ENTRY entrytime="00:01:07.00" eventid="1296" lane="2" heatid="8567" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNN" name="Cercle des Nageurs de Nyon" nation="SUI">
          <CONTACT city="Trelex" email="phil55@bluewin.ch" name="Mayer Philippe" phone="079 341 88 12" street="Chemin du treizou 7" zip="1270" />
          <ATHLETES>
            <ATHLETE birthdate="1955-01-01" firstname="Philippe" gender="M" lastname="Mayer" nation="SUI" license="4861" athleteid="7206">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="7347" lane="2" heatid="8592" />
                <ENTRY entrytime="NT" eventid="1196" lane="2" heatid="9736" />
                <ENTRY entrytime="00:02:46.18" eventid="1304" lane="5" heatid="8584" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOPR" name="Sport Figielski WOPR" nation="POL">
          <CONTACT country="PL" email="sport-figielski@02.pl" name="Grzegorz Figielski" />
          <ATHLETES>
            <ATHLETE birthdate="1958-01-01" firstname="Aleksandra" gender="F" lastname="Niespodziana" nation="POL" athleteid="7208">
              <ENTRIES>
                <ENTRY entrytime="00:02:55.00" eventid="1504" status="WDR" />
                <ENTRY entrytime="00:02:30.00" eventid="1054" status="WDR" />
                <ENTRY entrytime="00:00:35.00" eventid="1290" status="WDR" />
                <ENTRY entrytime="00:05:30.00" eventid="1072" status="WDR" />
                <ENTRY entrytime="00:01:20.00" eventid="1324" status="WDR" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Grzegorz" gender="M" lastname="Figielski" nation="POL" athleteid="7210">
              <ENTRIES>
                <ENTRY entrytime="00:03:00.00" eventid="1107" status="WDR" />
                <ENTRY entrytime="00:13:00.00" eventid="1196" status="WDR" />
                <ENTRY entrytime="00:06:00.00" eventid="1157" status="WDR" />
                <ENTRY entrytime="00:01:30.00" eventid="1342" status="WDR" />
                <ENTRY entrytime="00:03:20.00" eventid="1522" status="WDR" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="7211">
              <ENTRIES>
                <ENTRY entrytime="00:01:30.00" eventid="1342" lane="4" heatid="8600" />
                <ENTRY entrytime="NT" eventid="7347" lane="5" heatid="8592" />
                <ENTRY entrytime="00:02:50.00" eventid="1107" lane="3" heatid="8539" />
                <ENTRY entrytime="NT" eventid="1196" lane="4" heatid="9736" />
                <ENTRY entrytime="00:00:36.00" eventid="1292" lane="1" heatid="8559" />
                <ENTRY entrytime="00:00:31.00" eventid="1300" lane="2" heatid="8577" />
                <ENTRY entrytime="00:01:10.00" eventid="1450" status="DNS" lane="2" heatid="8622" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Jacek" gender="M" lastname="Adamski" nation="POL" athleteid="7212">
              <ENTRIES>
                <ENTRY entrytime="00:03:20.00" eventid="1522" status="WDR" />
                <ENTRY entrytime="00:01:30.00" eventid="1414" status="WDR" />
                <ENTRY entrytime="00:01:28.00" eventid="1296" status="WDR" />
                <ENTRY entrytime="00:03:35.00" eventid="1304" status="WDR" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1937-01-01" firstname="Zygmunt" gender="M" lastname="Lewandowski" nation="POL" athleteid="7213">
              <ENTRIES>
                <ENTRY entrytime="00:14:00.00" eventid="1196" status="WDR" />
                <ENTRY entrytime="00:03:40.00" eventid="1522" status="WDR" />
                <ENTRY entrytime="00:01:40.00" eventid="1342" status="WDR" />
                <ENTRY entrytime="00:01:40.00" eventid="1296" status="WDR" />
                <ENTRY entrytime="00:06:50.00" eventid="1157" status="WDR" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SVZ" name="Schwimmverein Zürileu" nation="SUI" region="RZO">
          <CONTACT city="Urdorf" email="billabongs@gmx.net" internet="www.svzuerileu.ch" name="Axel Mathis-Pairo" phone="+41 79 404 31 35" state="SUI" street="Untermatt 5" zip="8902" />
          <ATHLETES>
            <ATHLETE birthdate="1959-06-16" firstname="Heike" gender="F" lastname="Lischke" nation="GER" license="25770" athleteid="7288">
              <ENTRIES>
                <ENTRY entrytime="00:01:39.00" eventid="1396" lane="6" heatid="8611" />
                <ENTRY entrytime="00:01:26.60" eventid="1432" lane="3" heatid="8617" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SKL" name="Schwimmklub Luzern" nation="SUI">
          <CONTACT city="Horw" name="Krejci Josef" phone="041 340 33 42" street="Stegenstrasse 29" zip="6048" />
          <ATHLETES>
            <ATHLETE birthdate="1936-11-17" firstname="Olga" gender="F" lastname="Krejci" nation="SUI" license="2600" athleteid="7294">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.10" eventid="1298" lane="4" heatid="8571" />
                <ENTRY entrytime="00:00:52.50" eventid="1282" lane="2" heatid="8543" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1933-05-18" firstname="Josef" gender="M" lastname="Krejci" nation="SUI" license="5618" athleteid="7295">
              <ENTRIES>
                <ENTRY entrytime="00:03:10.00" eventid="1107" lane="3" heatid="8538" />
                <ENTRY entrytime="00:14:10.00" eventid="1196" lane="1" heatid="8589" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DUCKS" name="Duck&apos;s Creek" nation="RUS">
          <CONTACT email="info@dcsport.ru" name="Vera Tarasova" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Vladislav" gender="M" lastname="Bragin" nation="RUS" athleteid="7333">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.00" eventid="1296" lane="3" heatid="8567" />
                <ENTRY entrytime="00:00:28.20" eventid="1284" lane="3" heatid="8549" />
                <ENTRY entrytime="00:01:02.80" eventid="1414" status="DNS" lane="3" heatid="8615" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="POS" name="Poseydon" nation="RUS">
          <CONTACT email="info@dcsport.ru" name="Vera Tarasova" />
          <ATHLETES>
            <ATHLETE birthdate="1963-01-01" firstname="Vladislav" gender="M" lastname="Zagrebenko" nation="RUS" athleteid="7332">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.50" eventid="1284" lane="4" heatid="8549" />
                <ENTRY entrytime="00:01:09.50" eventid="1414" status="DNS" lane="2" heatid="8615" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-SSCHVB" name="Schweiz. Schwimmvereinigung" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1991-08-15" firstname="Michael" gender="M" lastname="Greber" nation="SUI" athleteid="7449">
              <HANDICAP breast="8" free="9" medley="9" />
              <ENTRIES>
                <ENTRY entrytime="00:01:02.63" eventid="1300" lane="1" heatid="8575" />
                <ENTRY entrytime="00:01:15.00" eventid="1378" lane="1" heatid="8606" />
                <ENTRY entrytime="00:02:23.13" eventid="1450" lane="2" heatid="8621" />
                <ENTRY entrytime="00:02:35.28" eventid="1288" lane="5" heatid="8554" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1964-11-01" firstname="Thomas" gender="M" lastname="Wittwer" nation="SUI" athleteid="7456">
              <HANDICAP breast="4" free="6" medley="6" />
              <ENTRIES>
                <ENTRY entrytime="00:01:02.00" eventid="1378" lane="5" heatid="8606" />
                <ENTRY entrytime="00:01:12.00" eventid="1284" lane="4" heatid="8545" />
                <ENTRY entrytime="00:02:05.00" eventid="1288" lane="2" heatid="8554" />
                <ENTRY entrytime="00:02:35.00" eventid="1414" lane="3" heatid="8612" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-30" firstname="Pablo" gender="M" lastname="Gallardo" nation="SUI" athleteid="7457">
              <HANDICAP free="9" />
              <ENTRIES>
                <ENTRY entrytime="00:06:58.00" eventid="1157" status="WDR" />
                <ENTRY entrytime="00:00:36.67" eventid="1300" status="WDR" />
                <ENTRY entrytime="00:01:25.00" eventid="1450" status="WDR" />
                <ENTRY entrytime="00:03:37.00" eventid="1107" status="WDR" />
                <ENTRY entrytime="00:14:22.00" eventid="1196" status="WDR" />
                <ENTRY entrytime="00:00:43.89" eventid="1292" status="WDR" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1959-08-31" firstname="Mirjam" gender="F" lastname="Schädler" nation="SUI" athleteid="7459">
              <HANDICAP free="6" />
              <ENTRIES>
                <ENTRY entrytime="00:04:46.00" eventid="1286" lane="2" heatid="8550" />
                <ENTRY entrytime="00:03:47.00" eventid="1432" lane="2" heatid="8616" />
                <ENTRY entrytime="00:01:42.00" eventid="1298" lane="3" heatid="8569" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-05-02" firstname="Dominik" gender="M" lastname="Stäger" nation="SUI" athleteid="7472">
              <HANDICAP breast="8" free="8" medley="8" />
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1107" lane="5" heatid="8538" />
                <ENTRY entrytime="NT" eventid="1378" lane="5" heatid="8605" />
                <ENTRY entrytime="NT" eventid="1288" lane="4" heatid="8553" />
                <ENTRY entrytime="NT" eventid="1450" lane="2" heatid="8620" />
                <ENTRY entrytime="NT" eventid="1300" lane="2" heatid="8574" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-13" firstname="Bruno" gender="M" lastname="Gasser" nation="SUI" athleteid="7475">
              <HANDICAP breast="10" free="10" medley="10" />
              <ENTRIES>
                <ENTRY entrytime="00:00:45.00" eventid="1300" lane="2" heatid="8575" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1961-02-05" firstname="Haenni" gender="M" lastname="Walter" nation="SUI" athleteid="7476">
              <HANDICAP breast="5" free="7" medley="6" />
              <ENTRIES>
                <ENTRY entrytime="00:02:28.00" eventid="1450" lane="5" heatid="8621" />
                <ENTRY entrytime="00:01:09.00" eventid="1300" lane="6" heatid="8575" />
                <ENTRY entrytime="00:01:12.00" eventid="1284" lane="2" heatid="8545" />
                <ENTRY entrytime="00:02:43.00" eventid="1414" lane="4" heatid="8612" />
                <ENTRY entrytime="00:01:25.00" eventid="1378" lane="3" heatid="8605" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1970-02-19" firstname="Denise" gender="F" lastname="Huser" nation="SUI" athleteid="7478">
              <HANDICAP breast="5" free="7" medley="7" />
              <ENTRIES>
                <ENTRY entrytime="00:03:18.00" eventid="1286" lane="3" heatid="8550" />
                <ENTRY entrytime="00:01:38.00" eventid="1360" lane="2" heatid="8603" />
                <ENTRY entrytime="00:01:44.00" eventid="1298" lane="4" heatid="8569" />
                <ENTRY entrytime="00:03:35.00" eventid="1432" lane="3" heatid="8616" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-14" firstname="Erwin" gender="M" lastname="Dürst" nation="SUI" athleteid="8527">
              <HANDICAP breast="8" free="9" medley="9" />
              <ENTRIES>
                <ENTRY entrytime="00:00:43.00" eventid="1300" lane="4" heatid="8575" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-WINT" name="Schwimmclub Winterthur Delfino" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1991-09-18" firstname="Stephanie" gender="F" lastname="Baumann" nation="SUI" athleteid="7450">
              <HANDICAP breast="9" free="9" medley="9" />
              <ENTRIES>
                <ENTRY entrytime="00:01:12.00" eventid="1432" lane="3" heatid="8618" />
                <ENTRY entrytime="00:00:33.00" eventid="1298" lane="3" heatid="8572" />
                <ENTRY entrytime="00:02:42.00" eventid="1054" lane="3" heatid="8536" />
                <ENTRY entrytime="00:01:28.00" eventid="1294" lane="3" heatid="8563" />
                <ENTRY entrytime="00:01:27.00" eventid="1286" lane="5" heatid="8552" />
                <ENTRY entrytime="00:03:06.00" eventid="1504" lane="4" heatid="8628" />
                <ENTRY entrytime="00:01:31.00" eventid="1324" lane="6" heatid="8599" />
                <ENTRY entrytime="00:05:40.00" eventid="1072" lane="3" heatid="8594" />
                <ENTRY entrytime="00:00:39.00" eventid="1360" lane="2" heatid="8604" />
                <ENTRY entrytime="00:01:42.00" eventid="1396" lane="3" heatid="8610" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-04-02" firstname="Lea" gender="F" lastname="Keller" nation="SUI" athleteid="7451">
              <HANDICAP breast="5" free="6" medley="6" />
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1054" lane="2" heatid="8535" />
                <ENTRY entrytime="00:03:41.00" eventid="1286" lane="4" heatid="8550" />
                <ENTRY entrytime="00:01:43.00" eventid="1282" lane="2" heatid="8542" />
                <ENTRY entrytime="00:01:46.00" eventid="1298" lane="2" heatid="8569" />
                <ENTRY entrytime="00:03:41.00" eventid="1396" lane="4" heatid="8609" />
                <ENTRY entrytime="00:03:45.00" eventid="1432" lane="4" heatid="8616" />
                <ENTRY entrytime="00:01:47.00" eventid="1360" lane="5" heatid="8603" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-10-18" firstname="Giuliana" gender="F" lastname="Bavaro" nation="SUI" athleteid="7452">
              <HANDICAP breast="7" free="8" />
              <ENTRIES>
                <ENTRY entrytime="00:01:19.00" eventid="1282" lane="3" heatid="8542" />
                <ENTRY entrytime="00:02:51.00" eventid="1396" lane="3" heatid="8609" />
                <ENTRY entrytime="00:01:58.00" eventid="1360" lane="1" heatid="8603" />
                <ENTRY entrytime="00:02:45.00" eventid="1432" lane="1" heatid="8617" />
                <ENTRY entrytime="00:01:28.00" eventid="1298" lane="6" heatid="8570" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-12-29" firstname="Ramona" gender="F" lastname="Loosli" nation="SUI" athleteid="7453">
              <HANDICAP breast="9" free="9" />
              <ENTRIES>
                <ENTRY entrytime="00:01:06.00" eventid="1282" lane="5" heatid="8543" />
                <ENTRY entrytime="00:02:03.00" eventid="1286" lane="2" heatid="8551" />
                <ENTRY entrytime="00:00:58.81" eventid="1360" lane="3" heatid="8603" />
                <ENTRY entrytime="00:02:17.00" eventid="1396" lane="5" heatid="8610" />
                <ENTRY entrytime="00:08:19.00" eventid="1072" lane="4" heatid="8593" />
                <ENTRY entrytime="00:00:50.68" eventid="1298" lane="6" heatid="8571" />
                <ENTRY entrytime="00:01:50.00" eventid="1432" lane="2" heatid="8617" />
                <ENTRY entrytime="NT" eventid="1294" lane="2" heatid="8562" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1991-07-14" firstname="Nicole" gender="F" lastname="Brunschwiler" nation="SUI" athleteid="7455">
              <HANDICAP breast="5" free="6" medley="6" />
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1282" lane="5" heatid="8542" />
                <ENTRY entrytime="NT" eventid="1360" lane="2" heatid="8602" />
                <ENTRY entrytime="NT" eventid="1286" lane="5" heatid="8550" />
                <ENTRY entrytime="NT" eventid="1298" lane="5" heatid="8569" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1990-12-04" firstname="Johannes" gender="M" lastname="Dumelin" nation="SUI" athleteid="7458">
              <HANDICAP breast="14" free="14" medley="14" />
              <ENTRIES>
                <ENTRY entrytime="00:01:25.00" eventid="1378" lane="4" heatid="8605" />
                <ENTRY entrytime="00:01:24.00" eventid="1284" lane="6" heatid="8545" />
                <ENTRY entrytime="00:03:13.00" eventid="1450" lane="3" heatid="8620" />
                <ENTRY entrytime="00:01:31.00" eventid="1300" lane="1" heatid="9290" />
                <ENTRY entrytime="NT" eventid="1414" lane="2" heatid="8612" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1987-12-15" firstname="Sabrina" gender="F" lastname="Pfeiffer" nation="SUI" athleteid="7462">
              <HANDICAP breast="201" free="201" medley="201" />
              <ENTRIES>
                <ENTRY entrytime="00:01:18.00" eventid="1298" lane="5" heatid="8570" />
                <ENTRY entrytime="00:01:08.00" eventid="1282" lane="1" heatid="8543" />
                <ENTRY entrytime="NT" eventid="1360" lane="4" heatid="8602" />
                <ENTRY entrytime="NT" eventid="1396" lane="2" heatid="8609" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-12-03" firstname="Carla" gender="F" lastname="De Bortoli" nation="SUI" athleteid="7468">
              <HANDICAP breast="13" free="13" medley="13" />
              <ENTRIES>
                <ENTRY entrytime="00:01:43.49" eventid="1396" lane="4" heatid="8610" />
                <ENTRY entrytime="00:00:48.53" eventid="1282" lane="6" heatid="8544" />
                <ENTRY entrytime="NT" eventid="1294" lane="4" heatid="8562" />
                <ENTRY entrytime="NT" eventid="1072" lane="2" heatid="8593" />
                <ENTRY entrytime="00:01:29.82" eventid="1432" lane="4" heatid="8617" />
                <ENTRY entrytime="00:00:40.79" eventid="1298" lane="2" heatid="8571" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-11-09" firstname="Nadin" gender="F" lastname="Lüthi" nation="SUI" athleteid="7471">
              <HANDICAP breast="9" free="9" medley="9" />
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1302" lane="1" heatid="8582" />
                <ENTRY entrytime="00:01:12.00" eventid="1282" lane="6" heatid="8543" />
                <ENTRY entrytime="00:02:23.00" eventid="1286" lane="1" heatid="8551" />
                <ENTRY entrytime="00:02:30.00" eventid="1396" lane="1" heatid="8610" />
                <ENTRY entrytime="00:01:20.00" eventid="1360" lane="4" heatid="8603" />
                <ENTRY entrytime="00:01:18.00" eventid="1298" lane="2" heatid="8570" />
                <ENTRY entrytime="00:02:12.00" eventid="1432" lane="5" heatid="8617" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1967-09-24" firstname="Wolf" gender="M" lastname="Schweitzer" nation="SUI" athleteid="7474">
              <HANDICAP breast="9" free="9" medley="9" />
              <ENTRIES>
                <ENTRY entrytime="00:02:58.00" eventid="1107" lane="2" heatid="8539" />
                <ENTRY entrytime="00:01:28.00" eventid="1414" lane="1" heatid="8614" />
                <ENTRY entrytime="00:00:31.00" eventid="1300" lane="4" heatid="8577" />
                <ENTRY entrytime="00:01:10.00" eventid="1450" lane="4" heatid="8622" />
                <ENTRY entrytime="NT" eventid="1292" lane="2" heatid="8558" />
                <ENTRY entrytime="00:00:41.90" eventid="1284" lane="2" heatid="8546" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-05" firstname="Philipp" gender="M" lastname="Rammerstorfer" nation="SUI" athleteid="7477">
              <HANDICAP breast="2" free="3" />
              <ENTRIES>
                <ENTRY entrytime="00:03:58.00" eventid="1288" lane="6" heatid="8554" />
                <ENTRY entrytime="00:01:36.00" eventid="1378" lane="2" heatid="8605" />
                <ENTRY entrytime="00:02:36.00" eventid="1284" lane="1" heatid="8545" />
                <ENTRY entrytime="00:03:52.00" eventid="1450" lane="4" heatid="8620" />
                <ENTRY entrytime="00:01:44.00" eventid="1300" lane="3" heatid="8574" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-CHUR" name="Schwimmclub Chur" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1994-04-26" firstname="Madlaina" gender="F" lastname="Gaudenz" nation="SUI" athleteid="7454">
              <HANDICAP breast="8" free="10" medley="9" />
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1290" lane="5" heatid="8557" />
                <ENTRY entrytime="NT" eventid="1294" lane="3" heatid="8562" />
                <ENTRY entrytime="00:01:32.00" eventid="1286" lane="6" heatid="8552" />
                <ENTRY entrytime="00:00:35.75" eventid="1298" lane="1" heatid="8572" />
                <ENTRY entrytime="00:01:19.00" eventid="1432" lane="1" heatid="8618" />
                <ENTRY entrytime="00:02:57.00" eventid="1054" lane="1" heatid="8536" />
                <ENTRY entrytime="00:06:00.00" eventid="1072" lane="5" heatid="8594" />
                <ENTRY entrytime="NT" eventid="1360" lane="3" heatid="8602" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-GER" name="Behindertenschwimmer Germany" nation="GER">
          <ATHLETES>
            <ATHLETE birthdate="1962-03-08" firstname="Markus" gender="M" lastname="Schnitzer" nation="GER" athleteid="7460">
              <HANDICAP free="10" medley="10" />
              <ENTRIES>
                <ENTRY entrytime="00:00:41.00" eventid="1378" lane="6" heatid="8607" />
                <ENTRY entrytime="00:02:50.00" eventid="1107" lane="4" heatid="8539" />
                <ENTRY entrytime="00:13:15.00" eventid="1196" lane="5" heatid="8589" />
                <ENTRY entrytime="00:06:20.00" eventid="1157" lane="4" heatid="8596" />
                <ENTRY entrytime="00:01:25.00" eventid="1288" lane="1" heatid="8555" />
                <ENTRY entrytime="00:01:35.00" eventid="1296" lane="5" heatid="8565" />
                <ENTRY entrytime="NT" eventid="1486" lane="2" heatid="8626" />
                <ENTRY entrytime="NT" eventid="1522" lane="6" heatid="8630" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-SKWORB" name="Schwimmklub Worb" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1978-02-12" firstname="Chantal" gender="F" lastname="Cavin" nation="SUI" athleteid="7461">
              <HANDICAP breast="11" free="11" medley="11" />
              <ENTRIES>
                <ENTRY entrytime="00:00:38.00" eventid="1290" lane="2" heatid="8557" />
                <ENTRY entrytime="00:01:30.00" eventid="1324" lane="1" heatid="8599" />
                <ENTRY entrytime="00:01:35.00" eventid="1294" lane="2" heatid="8563" />
                <ENTRY entrytime="00:00:45.00" eventid="1282" lane="1" heatid="8544" />
                <ENTRY entrytime="00:00:32.00" eventid="1298" lane="5" heatid="8573" />
                <ENTRY entrytime="00:01:11.00" eventid="1432" lane="6" heatid="8619" />
                <ENTRY entrytime="00:02:39.00" eventid="1054" lane="6" heatid="8537" />
                <ENTRY entrytime="00:05:50.00" eventid="1072" lane="2" heatid="8594" />
                <ENTRY entrytime="00:01:39.00" eventid="1396" status="WDR" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-SVK" name="Schwimmverein Kriens" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1990-05-08" firstname="Andrea" gender="F" lastname="Seiler" nation="SUI" athleteid="7463">
              <HANDICAP breast="9" free="9" medley="9" />
              <ENTRIES>
                <ENTRY entrytime="00:01:20.00" eventid="1432" lane="6" heatid="8618" />
                <ENTRY entrytime="00:00:41.00" eventid="1360" lane="1" heatid="8604" />
                <ENTRY entrytime="00:01:31.00" eventid="1286" lane="1" heatid="8552" />
                <ENTRY entrytime="00:03:23.00" eventid="1468" lane="2" heatid="8625" />
                <ENTRY entrytime="00:01:39.00" eventid="1294" lane="1" heatid="8563" />
                <ENTRY entrytime="00:00:35.00" eventid="1298" lane="5" heatid="8572" />
                <ENTRY entrytime="00:03:04.00" eventid="1054" lane="6" heatid="8536" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-BSGZ" name="Behindertensportgruppe Zimmerberg" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1984-11-23" firstname="Philipp" gender="M" lastname="Leuzinger" nation="SUI" athleteid="7464">
              <HANDICAP breast="9" free="9" medley="9" />
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1107" lane="4" heatid="8538" />
                <ENTRY entrytime="00:00:58.00" eventid="1300" lane="5" heatid="8575" />
                <ENTRY entrytime="NT" eventid="1288" lane="2" heatid="8553" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1983-08-07" firstname="Matthias" gender="M" lastname="Rusterholz" nation="SUI" athleteid="7465">
              <HANDICAP breast="9" free="9" medley="9" />
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1288" lane="3" heatid="8553" />
                <ENTRY entrytime="NT" eventid="1300" lane="6" heatid="8574" />
                <ENTRY entrytime="NT" eventid="1296" status="WDR" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1988-02-08" firstname="Nicole" gender="F" lastname="Odermatt" nation="SUI" athleteid="7466">
              <HANDICAP breast="7" free="7" medley="7" />
              <ENTRIES>
                <ENTRY entrytime="00:02:15.00" eventid="1286" lane="5" heatid="8551" />
                <ENTRY entrytime="00:00:58.00" eventid="1298" lane="3" heatid="8570" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1985-12-02" firstname="Cécile" gender="F" lastname="Bucher" nation="SUI" athleteid="7467">
              <HANDICAP breast="7" free="8" medley="8" />
              <ENTRIES>
                <ENTRY entrytime="00:02:25.00" eventid="1286" lane="6" heatid="8551" />
                <ENTRY entrytime="00:01:21.00" eventid="1298" lane="1" heatid="8570" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Basil" gender="M" lastname="Dias" nation="SUI" athleteid="7469">
              <HANDICAP breast="6" free="7" medley="7" />
              <ENTRIES>
                <ENTRY entrytime="00:02:19.00" eventid="1300" lane="4" heatid="8574" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1994-10-25" firstname="Svonislav" gender="M" lastname="Jankovic" nation="SUI" athleteid="7470">
              <HANDICAP breast="201" free="201" medley="201" />
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1300" lane="5" heatid="8574" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-LIMM" name="SV Limmat Sharks" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1974-07-03" firstname="Reto" gender="M" lastname="Thurnherr" nation="SUI" athleteid="7473">
              <HANDICAP breast="8" free="8" medley="8" />
              <ENTRIES>
                <ENTRY entrytime="00:06:00.00" eventid="1157" lane="5" heatid="8597" />
                <ENTRY entrytime="00:01:20.00" eventid="1450" lane="6" heatid="8622" />
                <ENTRY entrytime="00:00:40.00" eventid="1292" lane="3" heatid="8558" />
                <ENTRY entrytime="00:03:00.00" eventid="1107" lane="6" heatid="8539" />
                <ENTRY entrytime="00:00:36.00" eventid="1300" lane="1" heatid="8576" />
                <ENTRY entrytime="00:01:44.00" eventid="1296" lane="6" heatid="8565" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="H-BSGO" name="BSG Obwalden" nation="SUI">
          <ATHLETES>
            <ATHLETE birthdate="1985-08-17" firstname="Corinne" gender="F" lastname="Gasser" nation="SUI" athleteid="7479">
              <HANDICAP breast="14" free="14" medley="14" />
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="1298" lane="4" heatid="8570" />
                <ENTRY entrytime="00:01:30.00" eventid="1282" lane="4" heatid="8542" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SSG" name="SSG Saar MR" nation="GER">
          <CONTACT city="Friedrichsthal" country="DE" email="AnneSchmitt-SSG@web.de" name="Anne Schmitt" phone="0171 15 74 103" street="Ludwigstrasse 10" zip="66299" />
          <ATHLETES>
            <ATHLETE birthdate="1940-01-01" firstname="Hermann" gender="M" lastname="Sittner" nation="GER" license="93461" athleteid="7665">
              <ENTRIES>
                <ENTRY entrytime="00:04:18.00" eventid="1304" lane="5" heatid="8583" />
                <ENTRY entrytime="00:00:50.00" eventid="1284" lane="3" heatid="8545" />
                <ENTRY entrytime="00:01:55.00" eventid="1414" lane="5" heatid="8613" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TV 1872" name="TV 1872 Saarlouis" nation="FRA">
          <CONTACT city="Creutzwald" country="FR" name="Kurt Mayer" street="60 rue du Maréchal Ney" zip="57150" />
          <ATHLETES>
            <ATHLETE birthdate="1927-01-01" firstname="Kurt" gender="M" lastname="Mayer" nation="FRA" license="135080" athleteid="7670">
              <ENTRIES>
                <ENTRY entrytime="00:01:18.00" eventid="1378" lane="6" heatid="8606" />
                <ENTRY entrytime="00:06:12.00" eventid="1486" lane="4" heatid="8626" />
                <ENTRY entrytime="00:01:19.00" eventid="1284" lane="5" heatid="8545" />
                <ENTRY entrytime="00:02:54.00" eventid="1288" lane="1" heatid="8554" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GEN" name="Genève Natation 1885" nation="SUI" region="RSR">
          <CONTACT city="Genève 26" email="info@geneve-natation-1885.ch" fax="022/301.36.96" name="Secrétariat" phone="022/342.19.72" street="Piscine des Vernets" street2="Velardo Patricia" zip="CH-1211" />
          <ATHLETES>
            <ATHLETE birthdate="1959-07-18" firstname="Robert" gender="M" lastname="Alderton" nation="GBR" athleteid="7812">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.50" eventid="1378" status="DNS" lane="4" heatid="8608" />
                <ENTRY entrytime="00:01:10.00" eventid="1296" status="DNS" lane="3" heatid="8566" />
                <ENTRY entrytime="00:02:35.00" eventid="1486" status="DNS" lane="4" heatid="8627" />
                <ENTRY entrytime="00:00:35.00" eventid="1284" status="DNS" lane="5" heatid="8548" />
                <ENTRY entrytime="00:01:00.00" eventid="1288" status="DNS" lane="3" heatid="8556" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1970-12-12" firstname="Jonathan" gender="M" lastname="Banville" nation="CAN" license="15297" athleteid="7818">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.09" eventid="1414" lane="4" heatid="8615" />
                <ENTRY entrytime="00:02:20.09" eventid="1522" lane="3" heatid="8631" />
                <ENTRY entrytime="00:02:29.41" eventid="1304" lane="3" heatid="8584" />
                <ENTRY entrytime="00:01:03.29" eventid="1296" lane="4" heatid="8567" />
                <ENTRY entrytime="00:00:31.42" eventid="1284" lane="2" heatid="8549" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1975-08-06" firstname="Andreas" gender="M" lastname="Herty" nation="GER" license="18212" athleteid="7836">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.71" eventid="1378" lane="5" heatid="8608">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.80" eventid="1486" lane="6" heatid="8627">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.70" eventid="1296" lane="4" heatid="8566" />
                <ENTRY entrytime="00:01:14.20" eventid="1288" lane="5" heatid="8556" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-19" firstname="Daniela" gender="F" lastname="Menegon" nation="ITA" license="22084" athleteid="7847">
              <ENTRIES>
                <ENTRY entrytime="00:02:28.00" eventid="1054" lane="2" heatid="8537" />
                <ENTRY entrytime="00:00:31.60" eventid="1298" lane="2" heatid="8573" />
                <ENTRY entrytime="00:10:45.00" eventid="1177" lane="2" heatid="8588" />
                <ENTRY entrytime="00:05:15.00" eventid="1072" lane="5" heatid="8595" />
                <ENTRY entrytime="00:01:08.00" eventid="1432" lane="2" heatid="8619" />
                <ENTRY entrytime="00:03:00.00" eventid="1504" lane="3" heatid="8628" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1956-02-21" firstname="Simon" gender="M" lastname="Pagin" nation="SUI" license="16719" athleteid="7854">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.00" eventid="1284" lane="4" heatid="8546" />
                <ENTRY entrytime="00:01:26.00" eventid="1342" lane="3" heatid="8600" />
                <ENTRY entrytime="00:00:33.80" eventid="1292" lane="1" heatid="8560" />
                <ENTRY entrytime="00:00:31.00" eventid="1300" lane="3" heatid="8577" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="VN" name="Vevey Natation" nation="SUI">
          <CONTACT email="cmswisschris@gmail.com" name="Morgan Chris" />
          <ATHLETES>
            <ATHLETE birthdate="1969-01-01" firstname="Chris" gender="M" lastname="Morgan" nation="SUI" athleteid="7868">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.40" eventid="1292" lane="4" heatid="8561" />
                <ENTRY entrytime="00:00:26.70" eventid="1300" lane="5" heatid="8581" />
                <ENTRY entrytime="NT" eventid="1196" lane="6" heatid="8589" />
                <ENTRY entrytime="00:02:28.99" eventid="1107" lane="5" heatid="8540" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ASA" name="ASA Nuoto Cinisello ASD" nation="ITA">
          <CONTACT city="Cinisello Balsamo MI" country="IT" email="max.cassaghi@alice.it" name="Massimo Cassaghi" phone="0039 349 2259313" street="Via Vittorio Veneto 17" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Massimo" gender="M" lastname="Cassaghi" nation="ITA" license="LOM 035429" athleteid="7875">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.00" eventid="1378" lane="2" heatid="8608" />
                <ENTRY entrytime="00:00:59.50" eventid="1450" lane="5" heatid="8624" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOSIR" name="Mosir" nation="POL" shortname="MOSIR">
          <ATHLETES>
            <ATHLETE birthdate="1945-01-01" firstname="Jozef" gender="M" lastname="Rozalski" nation="POL" athleteid="7209">
              <ENTRIES>
                <ENTRY entrytime="00:03:45.00" eventid="1304" lane="4" heatid="8583" />
                <ENTRY entrytime="00:01:32.00" eventid="1342" lane="2" heatid="8600" />
                <ENTRY entrytime="00:01:35.00" eventid="1414" lane="6" heatid="8614" />
                <ENTRY entrytime="00:00:32.00" eventid="1300" lane="1" heatid="8577" />
                <ENTRY entrytime="00:03:25.00" eventid="1522" lane="1" heatid="8630" />
                <ENTRY entrytime="00:01:13.00" eventid="1450" lane="1" heatid="8622" />
                <ENTRY entrytime="00:01:24.00" eventid="1296" lane="6" heatid="8566" />
                <ENTRY entrytime="00:00:42.00" eventid="1284" lane="1" heatid="8546" />
                <ENTRY entrytime="00:00:34.00" eventid="1292" lane="3" heatid="8559" />
                <ENTRY entrytime="00:03:00.00" eventid="1107" lane="1" heatid="8539" />
                <ENTRY entrytime="00:06:20.00" eventid="1157" lane="2" heatid="8596" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="UNATTACHED" name="unattached">
          <OFFICIALS>
            <OFFICIAL officialid="7660" firstname="Christian" gender="M" grade="Schiiedsrichter A" lastname="Fahrni" />
          </OFFICIALS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
